netcdf clm_params_ed.c161103 {
dimensions:
	pft = 79 ;
	allpfts = 1 ;
	segment = 4 ;
	string_length = 40 ;
	variants = 2 ;
	litterclass = 6 ;
	param = 1 ;
	NCWD = 4 ;
variables:
	double FUN_fracfixers(pft) ;
	double Kmin_nh4(pft) ;
	double Kmin_no3(pft) ;
	double Vmax_nh4(pft) ;
	double Vmax_no3(pft) ;
	double a_fix(pft) ;
		a_fix:units = "unitless" ;
		a_fix:long_name = "An empirical curve-fitting parameter, which controls the shape of the symbiotic biological N fixation curve" ;
		a_fix:formula_terms = "Eq. (3) in Fisher et al (2010) and Eq.(5) in the Appendix of Brzostek et al (2014)" ;
		a_fix:references = "Houlton et al (2008); Fisher et al (2010); Brzostek et al (2014)" ;
	double aereoxid ;
		aereoxid:comment = "Use with the namelist switch use_aereoxid_prog.  If use_aereoxid_prog is equal to false, then read aereoxid from this parameter file.  Set to value between 0 & 1 (inclusive) for sensitivity tests." ;
		aereoxid:long_name = "Fraction of methane flux entering aerenchyma rhizosphere that will be oxidized rather than emitted" ;
		aereoxid:units = "unitless" ;
	double akc_active(pft) ;
		akc_active:units = "gC/m2" ;
		akc_active:long_name = "A parameter controls the cost as a function of root C (for the arbuscular mycorrhizal uptake pathway)" ;
		akc_active:formula_terms = "Eq. (3) and Table S2 from Brzostek et al (2014) and was tuned by M. Shi" ;
		akc_active:references = "Brzostek et al (2014)" ;
	double akn_active(pft) ;
		akn_active:units = "gN/m2" ;
		akn_active:long_name = "A parameter controls the cost as a function of soil N (for the arbuscular mycorrhizal uptake pathway)" ;
		akn_active:formula_terms = "Eq. (3) and Table S2 from Brzostek et al (2014) and was tuned by M. Shi" ;
		akn_active:references = "Brzostek et al (2014)" ;
	double aleaff(pft) ;
		aleaff:long_name = "Leaf Allocation coefficient parameter used in CNAllocationn" ;
		aleaff:units = "unitless" ;
		aleaff:coordinates = "pftname" ;
	double allconsl(pft) ;
		allconsl:long_name = "Leaf Allocation coefficient parameter power used in CNAllocation" ;
		allconsl:units = "unitless" ;
		allconsl:_FillValue = 0. ;
		allconsl:coordinates = "pftname" ;
	double allconss(pft) ;
		allconss:long_name = "Stem Allocation coefficient parameter power used in CNAllocation" ;
		allconss:units = "unitless" ;
		allconss:_FillValue = 0. ;
		allconss:coordinates = "pftname" ;
	double arootf(pft) ;
		arootf:long_name = "Root Allocation coefficient parameter used in CNAllocation" ;
		arootf:units = "unitless" ;
		arootf:_FillValue = 0. ;
		arootf:coordinates = "pftname" ;
	double arooti(pft) ;
		arooti:long_name = "Root Allocation coefficient parameter used in CNAllocation" ;
		arooti:units = "unitless" ;
		arooti:_FillValue = 0. ;
		arooti:coordinates = "pftname" ;
	double astemf(pft) ;
		astemf:long_name = "Stem Allocation coefficient parameter used in CNAllocation" ;
		astemf:units = "unitless" ;
		astemf:_FillValue = 0. ;
		astemf:coordinates = "pftname" ;
	double atmch4(allpfts) ;
		atmch4:long_name = "Atmospheric CH4 mixing ratio to prescribe if not provided by the atmospheric model" ;
		atmch4:units = "mol/mol" ;
	double b_fix(pft) ;
		b_fix:units = "unitless" ;
		b_fix:long_name = "An empirical curve-fitting parameter, which controls the shape of the symbiotic biological N fixation curve" ;
		b_fix:formula_terms = "Eq. (3) in Fisher et al (2010) and Eq.(5) in the Appendix of Brzostek et al (2014)" ;
		b_fix:references = "Houlton et al (2008); Fisher et al (2010); Brzostek et al (2014)" ;
	double baset(pft) ;
		baset:long_name = "Base Temperature, parameter used in accFlds" ;
		baset:units = "C" ;
		baset:coordinates = "pftname" ;
	double bdnr(allpfts) ;
		bdnr:long_name = "bulk denitrification rate" ;
		bdnr:units = "1/day" ;
	double bfact(pft) ;
		bfact:long_name = "Exponential factor used in CNAllocation for fraction allocated to leaf" ;
		bfact:units = "unitless" ;
		bfact:_FillValue = 0. ;
		bfact:coordinates = "pftname" ;
	double br_mr(allpfts) ;
		br_mr:long_name = "Base rate for maintenance respiration" ;
		br_mr:units = "gC/gN/s" ;
	double c3psn(pft) ;
		c3psn:long_name = "Photosynthetic pathway" ;
		c3psn:units = "flag" ;
		c3psn:coordinates = "pftname" ;
		c3psn:valid_range = 0., 1. ;
		c3psn:flag_meanings = "C4 C3" ;
		c3psn:flag_values = 0., 1. ;
	double c_fix(pft) ;
		c_fix:units = "unitless" ;
		c_fix:long_name = "An empirical curve-fitting parameter, which controls the shape of the symbiotic biological N fixation curve" ;
		c_fix:formula_terms = "Eq. (3) in Fisher et al (2010) and Eq.(5) in the Appendix of Brzostek et al (2014)" ;
		c_fix:references = "Houlton et al (2008); Fisher et al (2010); Brzostek et al (2014)" ;
	double capthick(allpfts) ;
		capthick:long_name = "Minimum thickness before assuming h2osfc is impermeable" ;
		capthick:units = "mm" ;
	double cc_dstem(pft) ;
		cc_dstem:units = "0 to 1" ;
		cc_dstem:long_name = "Combustion completeness factor for dead stem" ;
		cc_dstem:_FillValue = -999.99 ;
	double cc_leaf(pft) ;
		cc_leaf:units = "0 to 1" ;
		cc_leaf:long_name = "Combustion completeness factor for leaf" ;
		cc_leaf:_FillValue = -999.99 ;
	double cc_lstem(pft) ;
		cc_lstem:units = "0 to 1" ;
		cc_lstem:long_name = "Combustion completeness factor for live stem" ;
		cc_lstem:_FillValue = -999.99 ;
	double cc_other(pft) ;
		cc_other:units = "0 to 1" ;
		cc_other:long_name = "Combustion completeness factor for other plant" ;
		cc_other:_FillValue = -999.99 ;
	double ck(segment, pft) ;
		ck:coordinates = "segment pftname" ;
		ck:units = "unitless" ;
		ck:long_name = "weibull curve shape parameter" ;
	double cn_s1(allpfts) ;
		cn_s1:long_name = "C:N for SOM pool 1" ;
		cn_s1:units = "gC/gN" ;
	double cn_s1_bgc(allpfts) ;
		cn_s1_bgc:long_name = "C:N for SOM 1" ;
		cn_s1_bgc:units = "unitless" ;
	double cn_s2(allpfts) ;
		cn_s2:long_name = "C:N for SOM pool 2" ;
		cn_s2:units = "gC/gN" ;
	double cn_s2_bgc(allpfts) ;
		cn_s2_bgc:long_name = "C:N for SOM pool 2" ;
		cn_s2_bgc:units = "gC/gN" ;
	double cn_s3(allpfts) ;
		cn_s3:long_name = "C:N for SOM pool 3" ;
		cn_s3:units = "gC/gN" ;
	double cn_s3_bgc(allpfts) ;
		cn_s3_bgc:long_name = "C:N for SOM pool 3" ;
		cn_s3_bgc:units = "gC/gN" ;
	double cn_s4(allpfts) ;
		cn_s4:long_name = "C:N for SOM pool 4" ;
		cn_s4:units = "gC/gN" ;
	double cnscalefactor(allpfts) ;
		cnscalefactor:long_name = "Scale factor on CN decomposition for assigning methane flux" ;
		cnscalefactor:units = "unitless" ;
	double compet_decomp_nh4(allpfts) ;
		compet_decomp_nh4:long_name = "Relative competitiveness of immobilizers for NH4" ;
		compet_decomp_nh4:units = "unitless" ;
	double compet_decomp_no3(allpfts) ;
		compet_decomp_no3:long_name = "Relative competitiveness of immobilizers for NO3" ;
		compet_decomp_no3:units = "unitless" ;
	double compet_denit(allpfts) ;
		compet_denit:long_name = "Relative competitiveness of denitrifiers for NO3" ;
		compet_denit:units = "unitless" ;
	double compet_nit(allpfts) ;
		compet_nit:long_name = "Relative competitiveness of nitrifiers for NH4" ;
		compet_nit:units = "unitless" ;
	double compet_plant_nh4(allpfts) ;
		compet_plant_nh4:long_name = "Relative compettiveness of plants for NH4" ;
		compet_plant_nh4:units = "unitless" ;
	double compet_plant_no3(allpfts) ;
		compet_plant_no3:long_name = "Relative compettiveness of plants for NO3" ;
		compet_plant_no3:units = "unitless" ;
	double crit_dayl(allpfts) ;
		crit_dayl:long_name = "Critical day length for senescence" ;
		crit_dayl:units = "seconds" ;
	double crit_offset_fdd(allpfts) ;
		crit_offset_fdd:long_name = "Critical number of freezing days to initiate offset" ;
		crit_offset_fdd:units = "days" ;
	double crit_offset_swi(allpfts) ;
		crit_offset_swi:long_name = "Critical number of water stress days to initiate offset" ;
		crit_offset_swi:units = "days" ;
	double crit_onset_fdd(allpfts) ;
		crit_onset_fdd:long_name = "Critical number of freezing days to set gdd counter" ;
		crit_onset_fdd:units = "days" ;
	double crit_onset_swi(allpfts) ;
		crit_onset_swi:long_name = "Critical number of days > soilpsi_on for onset" ;
		crit_onset_swi:units = "days" ;
	double croot_stem(pft) ;
		croot_stem:long_name = "Allocation parameter: new coarse root C per new stem C" ;
		croot_stem:units = "gC/gC" ;
		croot_stem:coordinates = "pftname" ;
	double crop(pft) ;
		crop:long_name = "Binary crop PFT flag:" ;
		crop:units = "logical flag" ;
		crop:coordinates = "pftname" ;
		crop:valid_range = 0., 1. ;
		crop:flag_values = 0., 1. ;
		crop:flag_meanings = "NOT_crop crop_PFT" ;
	double cryoturb_diffusion_k(allpfts) ;
		cryoturb_diffusion_k:long_name = "The cryoturbation diffusive constant for vertical mixing of SOM" ;
		cryoturb_diffusion_k:units = "m^2/sec" ;
	double cwd_fcel(allpfts) ;
		cwd_fcel:long_name = "Cellulose fraction for CWD" ;
		cwd_fcel:units = "unitless" ;
	double cwd_flig(allpfts) ;
		cwd_flig:long_name = "Lignin fraction of coarse woody debris" ;
		cwd_flig:units = "unitless" ;
	double dayscrecover(allpfts) ;
		dayscrecover:long_name = "days to recover negative cpool" ;
		dayscrecover:units = "unitless" ;
	double deadwdcn(pft) ;
		deadwdcn:long_name = "Dead wood (xylem and heartwood) C:N" ;
		deadwdcn:units = "gC/gN" ;
		deadwdcn:coordinates = "pftname" ;
	double declfact(pft) ;
		declfact:long_name = "Decline factor for gddmaturity used in CNAllocation" ;
		declfact:units = "unitless" ;
		declfact:_FillValue = 0. ;
		declfact:coordinates = "pftname" ;
	double decomp_depth_efolding(allpfts) ;
		decomp_depth_efolding:long_name = "e-folding depth for reduction in decomposition. Sset to large number for depth-independance" ;
		decomp_depth_efolding:units = "m" ;
	double depth_runoff_Nloss(allpfts) ;
		depth_runoff_Nloss:long_name = "Depth over which runoff mixes with soil water for N loss to runoff" ;
		depth_runoff_Nloss:units = "m" ;
	double displar(pft) ;
		displar:long_name = "Ratio of displacement height to canopy top height" ;
		displar:units = "unitless" ;
		displar:coordinates = "pftname" ;
	double dleaf(pft) ;
		dleaf:long_name = "Characteristic leaf dimension" ;
		dleaf:units = "m" ;
		dleaf:coordinates = "pftname" ;
	double dnp(allpfts) ;
		dnp:long_name = "Denitrification proportion" ;
		dnp:units = "unitless" ;
	double dsladlai(pft) ;
		dsladlai:long_name = "Through canopy, projected area basis: dSLA/dLAI" ;
		dsladlai:units = "m^2/gC" ;
		dsladlai:coordinates = "pftname" ;
	double ef_time(allpfts) ;
		ef_time:long_name = "e-folding time constant" ;
		ef_time:units = "years" ;
	double ekc_active(pft) ;
		ekc_active:units = "gC/m2" ;
		ekc_active:long_name = "A parameter controls the cost as a function of root C (for the ectomycorrhizal uptake pathway)" ;
		ekc_active:formula_terms = "Eq. (3) and Table S2 from Brzostek et al (2014) and was tuned by M. Shi" ;
		ekc_active:references = "Brzostek et al (2014)" ;
	double ekn_active(pft) ;
		ekn_active:units = "gN/m2" ;
		ekn_active:long_name = "A parameter controls the cost as a function of soil N (for the ectomycorrhizal uptake pathway)" ;
		ekn_active:formula_terms = "Eq. (3) and Table S2 from Brzostek et al (2014) and was tuned by M. Shi" ;
		ekn_active:references = "Brzostek et al (2014)" ;
	double evergreen(pft) ;
		evergreen:long_name = "Binary flag for evergreen leaf habit" ;
		evergreen:units = "logical flag" ;
		evergreen:coordinates = "pftname" ;
		evergreen:flag_meanings = "NON-evergreen evergreen" ;
		evergreen:flag_values = 0., 1. ;
	double f_ch4(allpfts) ;
		f_ch4:long_name = "Ratio of CH4 production to total C mineralization" ;
		f_ch4:units = "unitless" ;
	double f_sat(allpfts) ;
		f_sat:long_name = "Volumetric soil water defining top of water table or where production is allowed" ;
		f_sat:units = "unitless" ;
	double fcur(pft) ;
		fcur:long_name = "Allocation parameter: fraction of allocation that goes to currently displayed growth, remainder to storage" ;
		fcur:units = "fraction" ;
		fcur:coordinates = "pftname" ;
	double fcurdv(pft) ;
		fcurdv:long_name = "Alternate fcur for use with CNDV" ;
		fcurdv:units = "fraction" ;
		fcurdv:coordinates = "pftname" ;
	double fd_pft(pft) ;
		fd_pft:units = "hr" ;
		fd_pft:long_name = "Fire duration" ;
		fd_pft:_FillValue = -999.99 ;
	double manunitro(pft) ;
		manunitro:long_name = "Max fertilizer to be applied in total" ;
		manunitro:units = "kg N/m2" ;
		manunitro:coordinates = "pftname" ;
	double ffrootcn(pft) ;
		ffrootcn:long_name = "Fine root C:N during organ fill" ;
		ffrootcn:units = "gC/gN" ;
		ffrootcn:coordinates = "pftname" ;
	double fleafcn(pft) ;
		fleafcn:long_name = "Leaf C:N during organ fill" ;
		fleafcn:units = "gC/gN" ;
		fleafcn:coordinates = "pftname" ;
	double fleafi(pft) ;
		fleafi:long_name = "Leaf Allocation coefficient parameter fraction used in CNAllocation" ;
		fleafi:units = "unitless" ;
		fleafi:_FillValue = 0. ;
		fleafi:coordinates = "pftname" ;
	double flivewd(pft) ;
		flivewd:long_name = "Allocation parameter: fraction of new wood that is live (phloem and ray parenchyma)" ;
		flivewd:units = "fraction" ;
		flivewd:coordinates = "pftname" ;
	double flnr(pft) ;
		flnr:long_name = "Fraction of leaf N in Rubisco enzyme" ;
		flnr:units = "fraction" ;
		flnr:coordinates = "pftname" ;
	double fm_droot(pft) ;
		fm_droot:units = "0 to 1" ;
		fm_droot:long_name = "Fire-related mortality factor for dead roots" ;
		fm_droot:_FillValue = -999.99 ;
	double fm_dstem(pft) ;
		fm_dstem:units = "0 to 1" ;
		fm_dstem:long_name = "Fire-related mortality factor for dead stem" ;
		fm_dstem:_FillValue = -999.99 ;
	double fm_leaf(pft) ;
		fm_leaf:units = "0 to 1" ;
		fm_leaf:long_name = "Fire-related mortality factor for leaf" ;
		fm_leaf:_FillValue = -999.99 ;
	double fm_lroot(pft) ;
		fm_lroot:units = "0 to 1" ;
		fm_lroot:long_name = "Fire-related mortality factor for live roots" ;
		fm_lroot:_FillValue = -999.99 ;
	double fm_lstem(pft) ;
		fm_lstem:units = "0 to 1" ;
		fm_lstem:long_name = "Fire-related mortality factor for live stem" ;
		fm_lstem:_FillValue = -999.99 ;
	double fm_other(pft) ;
		fm_other:units = "0 to 1" ;
		fm_other:long_name = "Fire-related mortality factor for other plant" ;
		fm_other:_FillValue = -999.99 ;
	double fm_root(pft) ;
		fm_root:units = "0 to 1" ;
		fm_root:long_name = "Fire-related mortality factor for fine roots" ;
		fm_root:_FillValue = -999.99 ;
	double fnitr(pft) ;
		fnitr:long_name = "Foliage nitrogen limitation factor" ;
		fnitr:units = "unitless" ;
		fnitr:coordinates = "pftname" ;
	double fr_fcel(pft) ;
		fr_fcel:long_name = "Fine root litter cellulose fraction" ;
		fr_fcel:units = "fraction" ;
		fr_fcel:coordinates = "pftname" ;
	double fr_flab(pft) ;
		fr_flab:long_name = "Fine root litter labile fraction" ;
		fr_flab:units = "fraction" ;
		fr_flab:coordinates = "pftname" ;
	double fr_flig(pft) ;
		fr_flig:long_name = "Fine root litter lignin fraction" ;
		fr_flig:units = "fraction" ;
		fr_flig:coordinates = "pftname" ;
	double froot_leaf(pft) ;
		froot_leaf:long_name = "Allocation parameter: new fine root C per new leaf C" ;
		froot_leaf:units = "gC/gC" ;
		froot_leaf:coordinates = "pftname" ;
	double frootcn(pft) ;
		frootcn:long_name = "Fine root C:N" ;
		frootcn:units = "gC/gN" ;
		frootcn:coordinates = "pftname" ;
	double frootcn_max(pft) ;
	double frootcn_min(pft) ;
	double froz_q10(allpfts) ;
		froz_q10:long_name = "Separate q10 for frozen soil respiration rates" ;
		froz_q10:units = "unitless" ;
	double fsr_pft(pft) ;
		fsr_pft:units = "m/s" ;
		fsr_pft:long_name = "Fire spread rate" ;
		fsr_pft:_FillValue = -999.99 ;
	double fstemcn(pft) ;
		fstemcn:long_name = "Stem C:N during organ fill" ;
		fstemcn:units = "gC/gN" ;
		fstemcn:coordinates = "pftname" ;
	double fstor2tran(allpfts) ;
		fstor2tran:long_name = "Fraction of storage to move to transfer for each onset" ;
		fstor2tran:units = "unitless" ;
	double fun_cn_flex_a(pft) ;
	double fun_cn_flex_b(pft) ;
	double fun_cn_flex_c(pft) ;
	double gddfunc_p1(allpfts) ;
		gddfunc_p1:long_name = "Parameter 1 to calculate GDD threshold as fn of annual T" ;
		gddfunc_p1:units = "unitless" ;
	double gddfunc_p2(allpfts) ;
		gddfunc_p2:long_name = "Parameter 2 to calculate GDD threshold as fn of annual T" ;
		gddfunc_p2:units = "unitless" ;
	double gddmin(pft) ;
		gddmin:long_name = "Minimim growing degree days used in CNPhenology" ;
		gddmin:units = "unitless" ;
		gddmin:_FillValue = 0. ;
		gddmin:coordinates = "pftname" ;
	double graincn(pft) ;
		graincn:long_name = "Grain C:N" ;
		graincn:units = "gC/gN" ;
		graincn:_FillValue = 0. ;
		graincn:coordinates = "pftname" ;
	double grnfill(pft) ;
		grnfill:long_name = "Grain fill parameter used in CNPhenology" ;
		grnfill:units = "unitless" ;
		grnfill:_FillValue = 0. ;
		grnfill:coordinates = "pftname" ;
	double grperc(pft) ;
		grperc:long_name = "Growth respiration factor" ;
		grperc:units = "unitless" ;
		grperc:coordinates = "pftname" ;
	double grpnow(pft) ;
		grpnow:long_name = "Growth respiration factor" ;
		grpnow:units = "unitless" ;
		grpnow:coordinates = "pftname" ;
	double highlatfact(allpfts) ;
		highlatfact:long_name = "Multiple of qflxlagd for high latitudes" ;
		highlatfact:units = "unitless" ;
	double hybgdd(pft) ;
		hybgdd:long_name = "Growing Degree Days for maturity used in CNPhenology" ;
		hybgdd:units = "unitless" ;
		hybgdd:_FillValue = 0. ;
		hybgdd:coordinates = "pftname" ;
	double i_flnr(pft) ;
	double i_vc(pft) ;
	double i_vca(pft) ;
	double i_vcad(pft) ;
	double irrigated(pft) ;
		irrigated:long_name = "Binary Irrigated PFT flag" ;
		irrigated:units = "logical flag" ;
		irrigated:coordinates = "pftname" ;
		irrigated:valid_range = 0., 1. ;
		irrigated:flag_meanings = "NOT_irrigated irrigated" ;
		irrigated:flag_values = 0., 1. ;
	double k_frag(allpfts) ;
		k_frag:long_name = "Fragmentation rate for CWD" ;
		k_frag:units = "1/day" ;
	double k_l1(allpfts) ;
		k_l1:long_name = "Decomposition rate for litter 1" ;
		k_l1:units = "1/day" ;
	double k_l2(allpfts) ;
		k_l2:long_name = "Decomposition rate for litter 2" ;
		k_l2:units = "1/day" ;
	double k_l3(allpfts) ;
		k_l3:long_name = "Decomposition rate for litter 3" ;
		k_l3:units = "1/day" ;
	double k_m(allpfts) ;
		k_m:long_name = "Michaelis-Menten oxidation rate constant for CH4 concentration" ;
		k_m:units = "mol/m3-w" ;
	double k_m_o2(allpfts) ;
		k_m_o2:long_name = "Michaelis-Menten oxidation rate constant for O2 concentration" ;
		k_m_o2:units = "mol/m3-w" ;
	double k_m_unsat(allpfts) ;
		k_m_unsat:long_name = "Michaelis-Menten oxidation rate constant for CH4 concentration" ;
		k_m_unsat:units = "mol/m3-w" ;
	double k_mort(allpfts) ;
		k_mort:long_name = "Coefficient of growth efficiency in mortality equation" ;
		k_mort:units = "unitless" ;
	double k_nitr_max(allpfts) ;
		k_nitr_max:long_name = "Maximum nitrification rate constant" ;
		k_nitr_max:units = "1/sec" ;
	double k_s1(allpfts) ;
		k_s1:long_name = "Decomposition rate for SOM 1" ;
		k_s1:units = "1/day" ;
	double k_s2(allpfts) ;
		k_s2:long_name = "Decomposition rate for SOM 2" ;
		k_s2:units = "1/day" ;
	double k_s3(allpfts) ;
		k_s3:long_name = "Decomposition rate for SOM 3" ;
		k_s3:units = "1/day" ;
	double k_s4(allpfts) ;
		k_s4:long_name = "Decomposition rate for SOM 4" ;
		k_s4:units = "1/day" ;
	double kc_nonmyc(pft) ;
		kc_nonmyc:units = "gC/m2" ;
		kc_nonmyc:long_name = "A parameter controls the cost as a function of root C (for the nonmycorrhizal uptake pathway)" ;
		kc_nonmyc:formula_terms = "Eq. (3) and Table S2 from Brzostek et al (2014) and was tuned by M. Shi" ;
		kc_nonmyc:references = "Brzostek et al (2014)" ;
	double kmax(segment, pft) ;
		kmax:coordinates = "segment pftname" ;
		kmax:units = "mm h2o (transpired)/mm h2o (water potential gradient)/sec" ;
		kmax:long_name = "plant segment max conductance" ;
	double kn_nonmyc(pft) ;
		kn_nonmyc:units = "gN/m2" ;
		kn_nonmyc:long_name = "A parameter controls the cost as a function of soil N (for the nonmycorrhizal uptake pathway)" ;
		kn_nonmyc:formula_terms = "Eq. (3) and Table S2 from Brzostek et al (2014) and was tuned by M. Shi" ;
		kn_nonmyc:references = "Brzostek et al (2014)" ;
	double kr_resorb(pft) ;
		kr_resorb:units = "gC/m2" ;
		kr_resorb:long_name = "A parameter controls the cost of retranslocation" ;
		kr_resorb:formula_terms = "Eq. (5) in Fisher et al (2010) and Eq. (6) in the Appendix of Brzostek et al (2014); was tuned by M. Shi for different phenological types of CLM" ;
		kr_resorb:references = "Fisher et al (2010); Brzostek et al (2014)" ;
	double krmax(pft) ;
		krmax:coordinates = "pftname" ;
		krmax:units = "mm h2o (transpired)/mm h2o (water potential gradient)/sec" ;
		krmax:long_name = "root segment max conductance" ;
	double laimx(pft) ;
		laimx:long_name = "Maximum Leaf Area Index used in CNVegStructUpdate" ;
		laimx:units = "unitless" ;
		laimx:_FillValue = 0. ;
		laimx:coordinates = "pftname" ;
	double lake_decomp_fact(allpfts) ;
		lake_decomp_fact:long_name = "Base decomposition rate (1/s) at 25oC in lake" ;
		lake_decomp_fact:units = "1/s" ;
	double leaf_long(pft) ;
		leaf_long:long_name = "Leaf longevity" ;
		leaf_long:units = "years" ;
		leaf_long:coordinates = "pftname" ;
	double leafcn(pft) ;
		leafcn:long_name = "Leaf C:N" ;
		leafcn:units = "gC/gN" ;
		leafcn:coordinates = "pftname" ;
	double leafcn_max(pft) ;
	double leafcn_min(pft) ;
	double lf_fcel(pft) ;
		lf_fcel:long_name = "Leaf litter cellulose fraction" ;
		lf_fcel:units = "fraction" ;
		lf_fcel:coordinates = "pftname" ;
	double lf_flab(pft) ;
		lf_flab:long_name = "Leaf litter labile fraction" ;
		lf_flab:units = "fraction" ;
		lf_flab:coordinates = "pftname" ;
	double lf_flig(pft) ;
		lf_flig:long_name = "Leaf litter lignin fraction" ;
		lf_flig:units = "fraction" ;
		lf_flig:coordinates = "pftname" ;
	double lfemerg(pft) ;
		lfemerg:long_name = "Leaf emergence parameter used in CNPhenology" ;
		lfemerg:units = "unitless" ;
		lfemerg:_FillValue = 0. ;
		lfemerg:coordinates = "pftname" ;
	double lflitcn(pft) ;
		lflitcn:long_name = "Leaf litter C:N" ;
		lflitcn:units = "gC/gN" ;
		lflitcn:coordinates = "pftname" ;
	double lfr_cn(pft) ;
	double livewdcn(pft) ;
		livewdcn:long_name = "Live wood (phloem and ray parenchyma) C:N" ;
		livewdcn:units = "gC/gN" ;
		livewdcn:coordinates = "pftname" ;
	double livewdcn_max(pft) ;
	double livewdcn_min(pft) ;
	double lmr_intercept_atkin(pft) ;
		lmr_intercept_atkin:long_name = "Intercept in the calculation of the top of canopy leaf maintenance respiration base rate. Original values from Atkin et al. in prep 2016." ;
		lmr_intercept_atkin:units = "umol CO2/m**2/s" ;
		lmr_intercept_atkin:coordinates = "pftname" ;
	double lwtop_ann(allpfts) ;
		lwtop_ann:long_name = "Live wood turnover proportion" ;
		lwtop_ann:units = "unitless" ;
	int max_NH_planting_date(pft) ;
		max_NH_planting_date:_FillValue = 0 ;
		max_NH_planting_date:long_name = "Maximum planting date for the Northern Hemipsphere" ;
		max_NH_planting_date:units = "YYYYMMDD" ;
		max_NH_planting_date:coordinates = "pftname" ;
		max_NH_planting_date:comment = "Typical U.S. latest planting dates according to AgroIBIS: Maize May 10th; soybean Jun 20th; spring wheat mid-May; winter wheat early Nov." ;
	int max_SH_planting_date(pft) ;
		max_SH_planting_date:_FillValue = 0 ;
		max_SH_planting_date:long_name = "Maximum planting date for the Southern Hemipsphere" ;
		max_SH_planting_date:units = "YYYYMMDD" ;
		max_SH_planting_date:coordinates = "pftname" ;
		max_SH_planting_date:comment = "Same as max_NH_planting_date, but offset by six months" ;
	double max_altdepth_cryoturbation(allpfts) ;
		max_altdepth_cryoturbation:long_name = "Maximum active layer thickness for cryoturbation to occur" ;
		max_altdepth_cryoturbation:units = "m" ;
	double max_altmultiplier_cryoturb(allpfts) ;
		max_altmultiplier_cryoturb:long_name = "Ratio of the maximum extent of cryoturbation to the active layer thickness" ;
		max_altmultiplier_cryoturb:units = "unitless" ;
	double maxpsi_hr(allpfts) ;
		maxpsi_hr:long_name = "Maximum soil water potential for heterotrophic resp" ;
		maxpsi_hr:units = "MPa" ;
	double mbbopt(pft) ;
		mbbopt:long_name = "Ball-Berry slope of conductance-photosynthesis relationship, unstressed" ;
		mbbopt:units = "umol H2O/umol CO2" ;
		mbbopt:coordinates = "pftname" ;
	double me_herb(allpfts) ;
		me_herb:long_name = "Moisture of extinction for herbaceous PFTs (proportion)" ;
		me_herb:units = "unitless" ;
	double me_woody(allpfts) ;
		me_woody:long_name = "Moisture of extinction for woody PFTs (proportion)" ;
		me_woody:units = "unitless" ;
	int mergetoclmpft(pft) ;
		mergetoclmpft:_FillValue = 0 ;
		mergetoclmpft:long_name = "CLM pft to merge this pft to" ;
		mergetoclmpft:units = "index" ;
		mergetoclmpft:coordinates = "pftname" ;
	int min_NH_planting_date(pft) ;
		min_NH_planting_date:_FillValue = 0 ;
		min_NH_planting_date:long_name = "Minimum planting date for the Northern Hemipsphere" ;
		min_NH_planting_date:units = "YYYYMMDD" ;
		min_NH_planting_date:coordinates = "pftname" ;
		min_NH_planting_date:comment = "Typical U.S. earliest planting dates according to AgroIBIS: Maize Apr 10th; soybean May 15th; spring wheat early Apr; winter wheat Sep 1st" ;
	int min_SH_planting_date(pft) ;
		min_SH_planting_date:_FillValue = 0 ;
		min_SH_planting_date:long_name = "Minimum planting date for the Southern Hemipsphere" ;
		min_SH_planting_date:units = "YYYYMMDD" ;
		min_SH_planting_date:coordinates = "pftname" ;
		min_SH_planting_date:comment = "Same as min_NH_planting_date, but offset by six months" ;
	double min_planting_temp(pft) ;
		min_planting_temp:long_name = "Average 5 day daily minimum temperature needed for planting" ;
		min_planting_temp:units = "K" ;
		min_planting_temp:coordinates = "pftname" ;
		min_planting_temp:_FillValue = 1000. ;
		min_planting_temp:comment = "From AGROIBIS derived from EPIC model parameterizations" ;
	double minfuel(allpfts) ;
		minfuel:long_name = "Dead fuel threshold to carry a fire" ;
		minfuel:units = "gC/m2" ;
	double mino2lim ;
		mino2lim:long_name = "Minimum anaerobic decomposition rate as a fraction of potential aerobic rate" ;
		mino2lim:units = "unitless" ;
	double minpsi_hr(allpfts) ;
		minpsi_hr:long_name = "Minimum soil water potential for heterotrophic resp" ;
		minpsi_hr:units = "MPa" ;
	int mxmat(pft) ;
		mxmat:_FillValue = 0 ;
		mxmat:long_name = "Maximum number of days to maturity parameter in CNPhenology" ;
		mxmat:units = "days" ;
		mxmat:coordinates = "pftname" ;
	double mxtmp(pft) ;
		mxtmp:long_name = "Max Temperature, parameter used in accFlds" ;
		mxtmp:units = "C" ;
		mxtmp:_FillValue = 0. ;
	double ndays_off(allpfts) ;
		ndays_off:long_name = "Number of days to complete leaf offset" ;
		ndays_off:units = "days" ;
	double ndays_on(allpfts) ;
		ndays_on:long_name = "Number of days to complete leaf onset" ;
		ndays_on:units = "days" ;
	double nfr_cn(pft) ;
	double nongrassporosratio(allpfts) ;
		nongrassporosratio:long_name = "Ratio of root porosity in non-grass to grass, used for aerenchyma transport" ;
		nongrassporosratio:units = "unitless" ;
	double organic_max(allpfts) ;
		organic_max:long_name = "Organic matter content where soil is assumed to act like peat for diffusion" ;
		organic_max:units = "kg/m3" ;
	double oxinhib(allpfts) ;
		oxinhib:long_name = "Inhibition of methane production by oxygen" ;
		oxinhib:units = "m^3/mol" ;
	double pHmax(allpfts) ;
		pHmax:long_name = "Maximum pH for methane production" ;
		pHmax:units = "unitless" ;
	double pHmin(allpfts) ;
		pHmin:long_name = "Minimum pH for methane production" ;
		pHmin:units = "unitless" ;
	double pconv(pft) ;
		pconv:long_name = "Deadstem proportions to send to conversion flux" ;
		pconv:units = "fraction" ;
		pconv:coordinates = "pftname" ;
		pconv:valid_range = 0., 1. ;
		pconv:comment = "pconv+pprod10+pprod100 must sum to 1.0" ;
	double perecm(pft) ;
		perecm:units = "unitless" ;
		perecm:long_name = "The percentage of the ectomycorrhizal-assciated plant of each PFT" ;
		perecm:ormula_terms = "Table 2 from Shi et al (in prep)" ;
		perecm:references = "Read (1991); Allen et al (1995); Phillips et al (2013)" ;
	char pftname(pft, string_length) ;
		pftname:long_name = "Description of plant type" ;
		pftname:units = "unitless" ;
	short pftnum(pft) ;
		pftnum:long_name = "Plant Functional Type number" ;
		pftnum:units = "unitless" ;
		pftnum:coordinates = "pftname" ;
	double pftpar20(pft) ;
		pftpar20:long_name = "Tree maximum crown area" ;
		pftpar20:units = "m2" ;
		pftpar20:_FillValue = 9999.9 ;
		pftpar20:coordinates = "pftname" ;
	double pftpar28(pft) ;
		pftpar28:long_name = "Minimum coldest monthly mean temperature" ;
		pftpar28:units = "degrees_Celsius" ;
		pftpar28:_FillValue = 9999.9 ;
		pftpar28:coordinates = "pftname" ;
	double pftpar29(pft) ;
		pftpar29:long_name = "Maximum coldest monthly mean temperature" ;
		pftpar29:units = "degrees_Celsius" ;
		pftpar29:_FillValue = 1000. ;
		pftpar29:coordinates = "pftname" ;
	double pftpar30(pft) ;
		pftpar30:long_name = "Minimum growing degree days (>= 5 degree Celsius)" ;
		pftpar30:units = "degree_C_days" ;
		pftpar30:coordinates = "pftname" ;
	double pftpar31(pft) ;
		pftpar31:long_name = "Upper limit of temperature of the warmest month (twmax)" ;
		pftpar31:units = "degrees_Celsius" ;
		pftpar31:_FillValue = 1000. ;
		pftpar31:coordinates = "pftname" ;
	double planting_temp(pft) ;
		planting_temp:long_name = "Average 10 day temperature needed for planting" ;
		planting_temp:units = "K" ;
		planting_temp:coordinates = "pftname" ;
		planting_temp:_FillValue = 1000. ;
		planting_temp:comment = "From AGROIBIS derived from EPIC model parameterizations" ;
	double porosmin(allpfts) ;
		porosmin:long_name = "Minimum aerenchyma porosity" ;
		porosmin:units = "unitless" ;
	double pprod10(pft) ;
		pprod10:long_name = "Deadstem proportions to send to 10 year product pool" ;
		pprod10:units = "fraction" ;
		pprod10:coordinates = "pftname" ;
		pprod10:valid_range = 0., 1. ;
		pprod10:comment = "pconv+pprod10+pprod100 must sum to 1.0" ;
	double pprod100(pft) ;
		pprod100:long_name = "Deadstem proportions to send to 100 year product pool" ;
		pprod100:units = "fraction" ;
		pprod100:coordinates = "pftname" ;
		pprod100:valid_range = 0., 1. ;
		pprod100:comment = "pconv+pprod10+pprod100 must sum to 1.0" ;
	double pprodharv10(pft) ;
		pprodharv10:long_name = "Deadstem proportions to send to 10 year harvest pool" ;
		pprodharv10:units = "fraction" ;
		pprodharv10:coordinates = "pftname" ;
		pprodharv10:_FillValue = 0. ;
		pprodharv10:valid_range = 0., 1. ;
		pprodharv10:comment = "100 year harvest is one minus this value" ;
	double psi50(segment, pft) ;
		psi50:coordinates = "segment pftname" ;
		psi50:units = "mm" ;
		psi50:long_name = "water potential at 50% loss of conductance" ;
	double psi_soil_ref(pft) ;
		psi_soil_ref:coordinates = "pftname" ;
		psi_soil_ref:units = "mm" ;
		psi_soil_ref:long_name = "water potential for calculating unstressed reference hydraulic conductivity, i.e., the no-stress soil water potential, the shape of the vulnerability curve function is defined by min(hk / hk@psi_soil_ref, 1.)" ;
	double q10_ch4oxid(allpfts) ;
		q10_ch4oxid:long_name = "Q10 oxidation constant" ;
		q10_ch4oxid:units = "unitless" ;
	double q10_hr(allpfts) ;
		q10_hr:long_name = "Q10 for heterotrophic respiration" ;
		q10_hr:units = "unitless" ;
	double q10_mr(allpfts) ;
		q10_mr:long_name = "Q10 for maintenance respiration" ;
		q10_mr:units = "unitless" ;
	double q10ch4(allpfts) ;
		q10ch4:long_name = "Q10 for methane production" ;
		q10ch4:units = "unitless" ;
	double q10ch4base ;
		q10ch4base:long_name = "Temperature at which the effective f_ch4 actually equals the constant f_ch4" ;
	double q10lakebase(allpfts) ;
		q10lakebase:long_name = "Base temperature for lake CH4 production" ;
		q10lakebase:units = "K" ;
	double qflxlagd(allpfts) ;
		qflxlagd:long_name = "Days to lag time-lagged surface runoff (qflx_surf_lag) in the tropics" ;
		qflxlagd:units = "days" ;
	double r_mort(allpfts) ;
		r_mort:long_name = "Mortality rate" ;
		r_mort:units = "1/year" ;
	double rc_npool(allpfts) ;
		rc_npool:long_name = "resistance for uptake from plant n pool" ;
		rc_npool:units = "unitless" ;
	double redoxlag(allpfts) ;
		redoxlag:long_name = "Number of days to lag in the calculation of finundated_lag" ;
		redoxlag:units = "days" ;
	double redoxlag_vertical(allpfts) ;
		redoxlag_vertical:long_name = "Time lag (days) to inhibit production for newly unsaturated layers" ;
		redoxlag_vertical:units = "days" ;
	double rf_cwdl2_bgc(allpfts) ;
		rf_cwdl2_bgc:long_name = "respiration fraction from CWD to litter 2" ;
		rf_cwdl2_bgc:units = "unitless" ;
	double rf_cwdl3_bgc(allpfts) ;
		rf_cwdl3_bgc:long_name = "respiration fraction from CWD to litter 3" ;
		rf_cwdl3_bgc:units = "unitless" ;
	double rf_l1s1(allpfts) ;
		rf_l1s1:long_name = "Respiration fraction for litter 1 -> SOM 1" ;
		rf_l1s1:units = "unitless" ;
	double rf_l1s1_bgc(allpfts) ;
		rf_l1s1_bgc:long_name = "Respiration fraction for litter 1 -> SOM 1" ;
		rf_l1s1_bgc:units = "unitless" ;
	double rf_l2s1_bgc(allpfts) ;
		rf_l2s1_bgc:long_name = "respiration fraction litter 2 to SOM 1" ;
		rf_l2s1_bgc:units = "unitless" ;
	double rf_l2s2(allpfts) ;
		rf_l2s2:long_name = "Respiration fraction for litter 2 -> SOM 2" ;
		rf_l2s2:units = "unitless" ;
	double rf_l3s2_bgc(allpfts) ;
		rf_l3s2_bgc:long_name = "respiration fraction from litter 3 to SOM 2" ;
		rf_l3s2_bgc:units = "unitless" ;
	double rf_l3s3(allpfts) ;
		rf_l3s3:long_name = "Respiration fraction for litter 3 -> SOM 3" ;
		rf_l3s3:units = "unitless" ;
	double rf_s1s2(allpfts) ;
		rf_s1s2:long_name = "Respiration fraction for SOM 1 -> SOM 2" ;
		rf_s1s2:units = "unitless" ;
	double rf_s2s1_bgc(allpfts) ;
		rf_s2s1_bgc:long_name = "respiration fraction SOM 2 to SOM 1" ;
		rf_s2s1_bgc:units = "unitless" ;
	double rf_s2s3(allpfts) ;
		rf_s2s3:long_name = "Respiration fraction for SOM 2 -> SOM 3" ;
		rf_s2s3:units = "unitless" ;
	double rf_s2s3_bgc(allpfts) ;
		rf_s2s3_bgc:long_name = "Respiration fraction for SOM 2 -> SOM 3" ;
		rf_s2s3_bgc:units = "unitless" ;
	double rf_s3s1_bgc(allpfts) ;
		rf_s3s1_bgc:long_name = "respiration fraction SOM 3 to SOM 1" ;
		rf_s3s1_bgc:units = "unitless" ;
	double rf_s3s4(allpfts) ;
		rf_s3s4:long_name = "Respiration fraction for SOM 3 -> SOM 4" ;
		rf_s3s4:units = "unitless" ;
	double rholnir(pft) ;
		rholnir:long_name = "Leaf reflectance: near-IR" ;
		rholnir:units = "fraction" ;
		rholnir:coordinates = "pftname" ;
	double rholvis(pft) ;
		rholvis:long_name = "Leaf reflectance: visible" ;
		rholvis:units = "fraction" ;
		rholvis:coordinates = "pftname" ;
	double rhosnir(pft) ;
		rhosnir:long_name = "Stem reflectance: near-IR" ;
		rhosnir:units = "fraction" ;
		rhosnir:coordinates = "pftname" ;
	double rhosvis(pft) ;
		rhosvis:long_name = "Stem reflectance: visible" ;
		rhosvis:units = "fraction" ;
		rhosvis:coordinates = "pftname" ;
	double rij_kro_a(allpfts) ;
		rij_kro_a:long_name = "Best-fit parameter of simple-structure model (Arah and Vinten 1995)" ;
		rij_kro_a:units = "unitless" ;
	double rij_kro_alpha(allpfts) ;
		rij_kro_alpha:long_name = "Simple-structure model parameter (Arah and Vinten 1995)" ;
		rij_kro_alpha:units = "unitless" ;
	double rij_kro_beta(allpfts) ;
		rij_kro_beta:long_name = "Simple-structure model parameter (Arah and Vinten 1995)" ;
		rij_kro_beta:units = "unitless" ;
	double rij_kro_delta(allpfts) ;
		rij_kro_delta:long_name = "Simple-structure model parameter (Arah and Vinten 1995)" ;
		rij_kro_delta:units = "unitless" ;
	double rij_kro_gamma(allpfts) ;
		rij_kro_gamma:long_name = "Simple-structure model parameter (Arah and Vinten 1995)" ;
		rij_kro_gamma:units = "unitless" ;
	double rob(allpfts) ;
		rob:long_name = "Ratio of root length to vertical depth (root obliquity)" ;
		rob:units = "unitless" ;
	double root_dmx(pft) ;
		root_dmx:long_name = "maximum rooting depth of crops" ;
		root_dmx:units = "m" ;
	double roota_par(pft) ;
		roota_par:long_name = "CLM rooting distribution parameter" ;
		roota_par:units = "1/m" ;
		roota_par:coordinates = "pftname" ;
	double rootb_par(pft) ;
		rootb_par:long_name = "CLM rooting distribution parameter" ;
		rootb_par:units = "1/m" ;
		rootb_par:coordinates = "pftname" ;
	double rootlitfrac(allpfts) ;
		rootlitfrac:long_name = "Fraction of soil organic matter associated with roots" ;
		rootlitfrac:units = "unitless" ;
	double s_fix(pft) ;
		s_fix:units = "gC/gN" ;
		s_fix:long_name = "A parameter controls the amount of the symtiotic biologcial N fixation uptake" ;
		s_fix:formula_terms = "Eq. (3) in Fisher et al (2010) and Eq.(5) in the Appendix of Brzostek et al (2014); was -30 in Brzostek et al (2014) and tuned to -60 by M. Shi" ;
		s_fix:references = "Houlton et al (2008); Fisher et al (2010); Brzostek et al (2014)" ;
	double s_flnr(pft) ;
	double s_vc(pft) ;
	double s_vca(pft) ;
	double s_vcad(pft) ;
	double satpow(allpfts) ;
		satpow:long_name = "Exponent on watsat for saturated soil solute diffusion" ;
		satpow:units = "unitless" ;
	double scale_factor_aere(allpfts) ;
		scale_factor_aere:long_name = "Scale factor on the aerenchyma area for sensitivity tests" ;
		scale_factor_aere:units = "unitless" ;
	double scale_factor_gasdiff(allpfts) ;
		scale_factor_gasdiff:long_name = "Scale factor for gas diffusion" ;
		scale_factor_gasdiff:units = "unitless" ;
	double scale_factor_liqdiff(allpfts) ;
		scale_factor_liqdiff:long_name = "Scale factor for solute diffusion in liquid (water)" ;
		scale_factor_liqdiff:units = "unitless" ;
	double season_decid(pft) ;
		season_decid:long_name = "Binary flag for seasonal-deciduous leaf habit" ;
		season_decid:units = "logical flag" ;
		season_decid:coordinates = "pftname" ;
		season_decid:flag_meanings = "NOT seasonal-deciduous" ;
		season_decid:flag_values = 0., 1. ;
	char segment(segment, string_length) ;
		segment:units = "unitless" ;
		segment:long_name = "description of hydraulic segment" ;
	double sf_minn(allpfts) ;
		sf_minn:long_name = "Soluble fraction of mineral N" ;
		sf_minn:units = "unitless" ;
	double sf_no3(allpfts) ;
		sf_no3:long_name = "Soluble fraction of NO3" ;
		sf_no3:units = "unitless" ;
	double shape_fluxprof_param1(allpfts) ;
		shape_fluxprof_param1:long_name = "Shape parameter of advection/diffusion profile" ;
		shape_fluxprof_param1:units = "unitless" ;
	double slatop(pft) ;
		slatop:long_name = "Specific Leaf Area (SLA) at top of canopy, projected area basis" ;
		slatop:units = "m^2/gC" ;
		slatop:coordinates = "pftname" ;
	double smp_crit(allpfts) ;
		smp_crit:long_name = "Critical soil moisture potential to reduce oxidation (mm) due to dessication of methanotrophs above the water table" ;
		smp_crit:units = "mm" ;
	double smpsc(pft) ;
		smpsc:long_name = "Soil water potential at full stomatal closure" ;
		smpsc:units = "mm" ;
		smpsc:coordinates = "pftname" ;
	double smpso(pft) ;
		smpso:long_name = "Soil water potential at full stomatal opening" ;
		smpso:units = "mm" ;
		smpso:coordinates = "pftname" ;
	double soilpsi_off(allpfts) ;
		soilpsi_off:long_name = "Critical soil water potential for leaf offset" ;
		soilpsi_off:units = "MPa" ;
	double soilpsi_on(allpfts) ;
		soilpsi_on:long_name = "Critical soil water potential for leaf onset" ;
		soilpsi_on:units = "MPa" ;
	double som_diffus(allpfts) ;
		som_diffus:long_name = "Vertical soil organic matter diffusion coefficient for flat adv/diff profile " ;
		som_diffus:units = "m^2/sec" ;
	double stem_leaf(pft) ;
		stem_leaf:long_name = "Allocation parameter: new stem C per new leaf C (-1 means use dynamic stem allocation)" ;
		stem_leaf:units = "gC/gC" ;
		stem_leaf:coordinates = "pftname" ;
	double stress_decid(pft) ;
		stress_decid:long_name = "Binary flag for stress-deciduous leaf habit" ;
		stress_decid:units = "logical flag" ;
		stress_decid:coordinates = "pftname" ;
		stress_decid:valid_range = 0., 1. ;
		stress_decid:flag_values = 0., 1. ;
		stress_decid:flag_meanings = "NOT stress_decidious" ;
	double surface_tension_water(allpfts) ;
		surface_tension_water:long_name = "Surface tension of water (Arah and Vinten 1995)" ;
		surface_tension_water:units = "J/m^2" ;
	double tau_cwd(allpfts) ;
		tau_cwd:long_name = "Corrected fragmentation rate constant CWD" ;
		tau_cwd:units = "1/year" ;
	double tau_l1(allpfts) ;
		tau_l1:long_name = "Turnover time of  litter 1" ;
		tau_l1:units = "year" ;
	double tau_l2_l3(allpfts) ;
		tau_l2_l3:long_name = "Turnover time of  litter 2 and litter 3" ;
		tau_l2_l3:units = "year" ;
	double tau_s1(allpfts) ;
		tau_s1:long_name = "Turnover time of soil organic matter (SOM) 1" ;
		tau_s1:units = "year" ;
	double tau_s2(allpfts) ;
		tau_s2:long_name = "Turnover time of soil organic matter (SOM) 2" ;
		tau_s2:units = "year" ;
	double tau_s3(allpfts) ;
		tau_s3:long_name = "Turnover time of soil organic matter (SOM) 3" ;
		tau_s3:units = "year" ;
	double taulnir(pft) ;
		taulnir:long_name = "Leaf transmittance: near-IR" ;
		taulnir:units = "fraction" ;
		taulnir:coordinates = "pftname" ;
	double taulvis(pft) ;
		taulvis:long_name = "Leaf transmittance: visible" ;
		taulvis:units = "fraction" ;
		taulvis:coordinates = "pftname" ;
	double tausnir(pft) ;
		tausnir:long_name = "Stem transmittance: near-IR" ;
		tausnir:units = "fraction" ;
		tausnir:coordinates = "pftname" ;
	double tausvis(pft) ;
		tausvis:long_name = "Stem transmittance: visible" ;
		tausvis:units = "fraction" ;
		tausvis:coordinates = "pftname" ;
	double unsat_aere_ratio(allpfts) ;
		unsat_aere_ratio:long_name = "Ratio to multiply upland vegetation aerenchyma porosity by compared to inundated systems" ;
		unsat_aere_ratio:units = "unitless" ;
	double vgc_max(allpfts) ;
		vgc_max:long_name = "Ratio of saturation pressure triggering ebullition" ;
		vgc_max:units = "unitless" ;
	double vmax_ch4_oxid(allpfts) ;
		vmax_ch4_oxid:long_name = "Oxidation rate constant" ;
		vmax_ch4_oxid:units = "mol/m3-w/s" ;
	double vmax_oxid_unsat(allpfts) ;
		vmax_oxid_unsat:long_name = "Oxidation rate constant" ;
		vmax_oxid_unsat:units = "mol/m3-w/s" ;
	double wcf(allpfts) ;
		wcf:long_name = "Wood combustion fraction" ;
		wcf:units = "unitless" ;
	double woody(pft) ;
		woody:long_name = "Binary woody lifeform flag" ;
		woody:units = "logical flag" ;
		woody:coordinates = "pftname" ;
		woody:valid_range = 0., 1. ;
		woody:flag_values = 0., 1. ;
		woody:flag_meanings = "NON_woody woody" ;
	double xl(pft) ;
		xl:long_name = "Leaf/stem orientation index" ;
		xl:units = "unitless" ;
		xl:coordinates = "pftname" ;
		xl:valid_range = -1., 1. ;
	double z0mr(pft) ;
		z0mr:long_name = "Ratio of momentum roughness length to canopy top height" ;
		z0mr:units = "unitless" ;
		z0mr:coordinates = "pftname" ;
	double ztopmx(pft) ;
		ztopmx:long_name = "Canopy top coefficient used in CNVegStructUpdate" ;
		ztopmx:units = "m" ;
		ztopmx:_FillValue = 0. ;
		ztopmx:coordinates = "pftname" ;
	double rootprof_beta(variants, pft) ;
		rootprof_beta:long_name = "Rooting beta parameter, for C and N vertical discretization" ;
		rootprof_beta:units = "unitless" ;
	double wood_density(pft) ;
	double BB_slope(pft) ;
	double alpha_stem(pft) ;
	double leaf_stor_priority(pft) ;
	double max_dbh(pft) ;
	double cushion(pft) ;
	double hgt_min(pft) ;
	double freezetol(pft) ;
	double resp_drought_response(pft) ;
	double leafwatermax(pft) ;
	double rootresist(pft) ;
	double soilbeta(pft) ;
	double crown(pft) ;
	double bark_scaler(pft) ;
	double crown_kill(pft) ;
	double initd(pft) ;
	double sd_mort(pft) ;
	double seed_rain(pft) ;
	double bb_slope(pft) ;
	double root_long(pft) ;
	double seed_alloc(pft) ;
	double clone_alloc(pft) ;
	double sapwood_ratio(pft) ;
	double grass_spread(param) ;
	double comp_excln(param) ;
	double stress_mort(param) ;
	double dispersal(param) ;
	double gr_perc(param) ;
	double maxspread(param) ;
	double minspread(param) ;
	double init_litter(param) ;
	double nfires(param) ;
	double understorey_death(param) ;
	double profile_tol(param) ;
	double ag_biomass(param) ;
	double alpha_FMC(litterclass) ;
	double SAV(litterclass) ;
	double FBD(litterclass) ;
	double max_decomp(litterclass) ;
	double min_moisture(litterclass) ;
	double mid_moisture(litterclass) ;
	double low_moisture_C(litterclass) ;
	double low_moisture_S(litterclass) ;
	double mid_moisture_C(litterclass) ;
	double mid_moisture_S(litterclass) ;
	double CWD_frac(NCWD) ;
	double fdi_a ;
	double fdi_b ;
	double fdi_alpha ;
	double miner_total ;
	double fuel_energy ;
	double part_dens ;
	double miner_damp ;
	double max_durat ;
	double durat_slope ;
	double alpha_SH ;

// global attributes:
		:Conventions = "CF-1.0" ;
		:title = "Vegetation (Plant Function Type or PFT) constants" ;
		:nco_openmp_thread_number = 1 ;
		:history = "Thu Nov  3 15:34:37 2016: ncrename -v fertnitro,manunitro /glade/p/cesm/cseg/inputdata/lnd/clm2/paramdata/clm_params_ed.c160808.nc /glade/p/cesm/cseg/inputdata/lnd/clm2/paramdata/clm_params_ed.c161103.nc" ;
		:NCO = "\"4.5.5\"" ;
data:

 FUN_fracfixers = 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5 ;

 Kmin_nh4 = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Kmin_no3 = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Vmax_nh4 = 2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 
    2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 
    2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 
    2.7e-08, 2.7e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Vmax_no3 = 2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 
    2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 
    2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 2.7e-08, 
    2.7e-08, 2.7e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 a_fix = -3.61999988555908, -3.61999988555908, -3.61999988555908, 
    -3.61999988555908, -3.61999988555908, -3.61999988555908, 
    -3.61999988555908, -3.61999988555908, -3.61999988555908, 
    -3.61999988555908, -3.61999988555908, -3.61999988555908, 
    -3.61999988555908, -3.61999988555908, -3.61999988555908, 
    -3.61999988555908, -3.61999988555908, -3.61999988555908, 
    -3.61999988555908, -3.61999988555908, -3.61999988555908, 
    -3.61999988555908, -3.61999988555908, -3.61999988555908, 
    -3.61999988555908, -3.61999988555908, -3.61999988555908, 
    -3.61999988555908, -3.61999988555908, -3.61999988555908, 
    -3.61999988555908, -3.61999988555908, -3.61999988555908, 
    -3.61999988555908, -3.61999988555908, -3.61999988555908, 
    -3.61999988555908, -3.61999988555908, -3.61999988555908, 
    -3.61999988555908, -3.61999988555908, -3.61999988555908, 
    -3.61999988555908, -3.61999988555908, -3.61999988555908, 
    -3.61999988555908, -3.61999988555908, -3.61999988555908, 
    -3.61999988555908, -3.61999988555908, -3.61999988555908, 
    -3.61999988555908, -3.61999988555908, -3.61999988555908, 
    -3.61999988555908, -3.61999988555908, -3.61999988555908, 
    -3.61999988555908, -3.61999988555908, -3.61999988555908, 
    -3.61999988555908, -3.61999988555908, -3.61999988555908, 
    -3.61999988555908, -3.61999988555908, -3.61999988555908, 
    -3.61999988555908, -3.61999988555908, -3.61999988555908, 
    -3.61999988555908, -3.61999988555908, -3.61999988555908, 
    -3.61999988555908, -3.61999988555908, -3.61999988555908, 
    -3.61999988555908, -3.61999988555908, -3.61999988555908, -3.61999988555908 ;

 aereoxid = 0 ;

 akc_active = 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137, 0.000488954601190137, 
    0.000488954601190137, 0.000488954601190137 ;

 akn_active = 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589, 0.000438282092653589, 
    0.000438282092653589, 0.000438282092653589 ;

 aleaff = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 allconsl = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 5, 5, 3, 3, 3, 
    3, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, 2, 2, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 3, 3, _, _, _, _, 5, 5, _, 
    _, _, _, _, _, 5, 5, 2, 2 ;

 allconss = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 1, 1, 1, 
    1, 5, 5, 1, 1, 1, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, 5, 5, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 1, 1, _, _, _, _, 2, 2, _, 
    _, _, _, _, _, 2, 2, 5, 5 ;

 arootf = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0.05, 0.05, _, 
    _, _, _, 0.2, 0.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0.2, 
    0.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, 0.05, 0.05, _, _, _, _, _, _, 0.05, 0.05, 0.2, 0.2 ;

 arooti = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0.4, 0.4, 0.3, 
    0.3, 0.3, 0.3, 0.5, 0.5, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, _, _, _, 
    _, _, _, _, _, 0.5, 0.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, 0.3, 0.3, _, _, _, _, 0.4, 0.4, _, _, _, _, _, _, 0.4, 0.4, 0.5, 0.5 ;

 astemf = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0.05, 
    0.05, 0.05, 0.05, 0.3, 0.3, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, _, _, _, _, _, _, _, _, 0.3, 0.3, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, 0.05, 0.05, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, 0.3, 0.3 ;

 atmch4 = 1.7e-06 ;

 b_fix = 0.270000010728836, 0.270000010728836, 0.270000010728836, 
    0.270000010728836, 0.270000010728836, 0.270000010728836, 
    0.270000010728836, 0.270000010728836, 0.270000010728836, 
    0.270000010728836, 0.270000010728836, 0.270000010728836, 
    0.270000010728836, 0.270000010728836, 0.270000010728836, 
    0.270000010728836, 0.270000010728836, 0.270000010728836, 
    0.270000010728836, 0.270000010728836, 0.270000010728836, 
    0.270000010728836, 0.270000010728836, 0.270000010728836, 
    0.270000010728836, 0.270000010728836, 0.270000010728836, 
    0.270000010728836, 0.270000010728836, 0.270000010728836, 
    0.270000010728836, 0.270000010728836, 0.270000010728836, 
    0.270000010728836, 0.270000010728836, 0.270000010728836, 
    0.270000010728836, 0.270000010728836, 0.270000010728836, 
    0.270000010728836, 0.270000010728836, 0.270000010728836, 
    0.270000010728836, 0.270000010728836, 0.270000010728836, 
    0.270000010728836, 0.270000010728836, 0.270000010728836, 
    0.270000010728836, 0.270000010728836, 0.270000010728836, 
    0.270000010728836, 0.270000010728836, 0.270000010728836, 
    0.270000010728836, 0.270000010728836, 0.270000010728836, 
    0.270000010728836, 0.270000010728836, 0.270000010728836, 
    0.270000010728836, 0.270000010728836, 0.270000010728836, 
    0.270000010728836, 0.270000010728836, 0.270000010728836, 
    0.270000010728836, 0.270000010728836, 0.270000010728836, 
    0.270000010728836, 0.270000010728836, 0.270000010728836, 
    0.270000010728836, 0.270000010728836, 0.270000010728836, 
    0.270000010728836, 0.270000010728836, 0.270000010728836, 0.270000010728836 ;

 baset = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 8, 0, 0, 0, 0, 
    10, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 10, 0, 0, 0, 0, 10, 10, 
    0, 0, 0, 0, 0, 0, 10, 10, 10, 10 ;

 bdnr = 0.5 ;

 bfact = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0.1, 0.1, 0.1, 
    0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 
    0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 
    0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 
    0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 
    0.1, 0.1, 0.1 ;

 br_mr = 2.525e-06 ;

 c3psn = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 0, 0, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 1, 1, 
    1, 1, 1, 1, 0, 0, 1, 1 ;

 c_fix = 25.1499996185303, 25.1499996185303, 25.1499996185303, 
    25.1499996185303, 25.1499996185303, 25.1499996185303, 25.1499996185303, 
    25.1499996185303, 25.1499996185303, 25.1499996185303, 25.1499996185303, 
    25.1499996185303, 25.1499996185303, 25.1499996185303, 25.1499996185303, 
    25.1499996185303, 25.1499996185303, 25.1499996185303, 25.1499996185303, 
    25.1499996185303, 25.1499996185303, 25.1499996185303, 25.1499996185303, 
    25.1499996185303, 25.1499996185303, 25.1499996185303, 25.1499996185303, 
    25.1499996185303, 25.1499996185303, 25.1499996185303, 25.1499996185303, 
    25.1499996185303, 25.1499996185303, 25.1499996185303, 25.1499996185303, 
    25.1499996185303, 25.1499996185303, 25.1499996185303, 25.1499996185303, 
    25.1499996185303, 25.1499996185303, 25.1499996185303, 25.1499996185303, 
    25.1499996185303, 25.1499996185303, 25.1499996185303, 25.1499996185303, 
    25.1499996185303, 25.1499996185303, 25.1499996185303, 25.1499996185303, 
    25.1499996185303, 25.1499996185303, 25.1499996185303, 25.1499996185303, 
    25.1499996185303, 25.1499996185303, 25.1499996185303, 25.1499996185303, 
    25.1499996185303, 25.1499996185303, 25.1499996185303, 25.1499996185303, 
    25.1499996185303, 25.1499996185303, 25.1499996185303, 25.1499996185303, 
    25.1499996185303, 25.1499996185303, 25.1499996185303, 25.1499996185303, 
    25.1499996185303, 25.1499996185303, 25.1499996185303, 25.1499996185303, 
    25.1499996185303, 25.1499996185303, 25.1499996185303, 25.1499996185303 ;

 capthick = 100 ;

 cc_dstem = 0, 0.22, 0.25, 0.25, 0.22, 0.22, 0.22, 0.22, 0.22, 0.3, 0.3, 0.3, 
    0.8, 0.8, 0.8, 0.8, 0.8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 cc_leaf = 0, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 
    0.8, 0.8, 0.8, 0.8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 cc_lstem = 0, 0.22, 0.25, 0.25, 0.22, 0.22, 0.22, 0.22, 0.22, 0.3, 0.3, 0.3, 
    0.8, 0.8, 0.8, 0.8, 0.8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 cc_other = 0, 0.45, 0.5, 0.5, 0.45, 0.45, 0.45, 0.45, 0.45, 0.55, 0.55, 
    0.55, 0.8, 0.8, 0.8, 0.8, 0.8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ck =
  0, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 
    3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 
    3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 
    3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 
    3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 
    3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 
    3.95, 3.95, 3.95, 3.95, 3.95, 3.95,
  0, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 
    3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 
    3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 
    3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 
    3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 
    3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 
    3.95, 3.95, 3.95, 3.95, 3.95, 3.95,
  0, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 
    3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 
    3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 
    3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 
    3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 
    3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 
    3.95, 3.95, 3.95, 3.95, 3.95, 3.95,
  0, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 
    3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 
    3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 
    3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 
    3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 
    3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 3.95, 
    3.95, 3.95, 3.95, 3.95, 3.95, 3.95 ;

 cn_s1 = 12 ;

 cn_s1_bgc = 8 ;

 cn_s2 = 12 ;

 cn_s2_bgc = 11 ;

 cn_s3 = 10 ;

 cn_s3_bgc = 11 ;

 cn_s4 = 10 ;

 cnscalefactor = 1 ;

 compet_decomp_nh4 = 1 ;

 compet_decomp_no3 = 1 ;

 compet_denit = 1 ;

 compet_nit = 1 ;

 compet_plant_nh4 = 1 ;

 compet_plant_no3 = 1 ;

 crit_dayl = 39300 ;

 crit_offset_fdd = 15 ;

 crit_offset_swi = 15 ;

 crit_onset_fdd = 15 ;

 crit_onset_swi = 15 ;

 croot_stem = 0, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 crop = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1 ;

 cryoturb_diffusion_k = 1.5855e-11 ;

 cwd_fcel = 0.76 ;

 cwd_flig = 0.24 ;

 dayscrecover = 30 ;

 deadwdcn = 1, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 0, 0, 
    0, 0, 0, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 
    500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 
    500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 
    500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 500, 
    500, 500, 500, 500, 500, 500, 500 ;

 declfact = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 1.05, 1.05, 
    1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 
    1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 
    1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 
    1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 
    1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05, 1.05 ;

 decomp_depth_efolding = 0.5 ;

 depth_runoff_Nloss = 0.05 ;

 displar = 0, 0.67, 0.67, 0.67, 0.67, 0.67, 0.67, 0.67, 0.67, 0.68, 0.68, 
    0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 
    0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 
    0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 
    0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 
    0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 
    0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68, 0.68 ;

 dleaf = 0, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 
    0.04, 0.04, 0.04, 0.04, 0.04, 0.04, 0.04 ;

 dnp = 0.01 ;

 dsladlai = 0, 0.00125, 0.001, 0.003, 0.0015, 0.0015, 0.004, 0.004, 0.004, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ef_time = 1 ;

 ekc_active = 0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806, 0.0104575719776806, 0.0104575719776806, 
    0.0104575719776806 ;

 ekn_active = 0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583, 0.00183577041869583, 0.00183577041869583, 
    0.00183577041869583 ;

 evergreen = 0, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 f_ch4 = 0.2 ;

 f_sat = 0.95 ;

 fcur = 0, 1, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1 ;

 fcurdv = 0, 1, 1, 0.5, 1, 1, 0.5, 0.5, 0.5, 1, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 fd_pft = 0, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 manunitro = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0149999996647239, 0.0149999996647239, 0.00800000037997961, 
    0.00800000037997961, 0.00800000037997961, 0.00800000037997961, 
    0.00249999994412065, 0.00249999994412065, 0.00800000037997961, 
    0.00800000037997961, 0.00800000037997961, 0.00800000037997961, 
    0.00800000037997961, 0.00800000037997961, 0.00800000037997961, 
    0.00800000037997961, 0, 0, 0, 0, 0, 0, 0, 0, 0.02, 0.02, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02, 0.02, 0, 0, 0, 0, 0.04, 
    0.04, 0, 0, 0, 0, 0, 0, 0.03, 0.03, 0.05, 0.05 ;

 ffrootcn = 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 
    999, 999, 999, 999, 0, 0, 40, 40, 40, 40, 0, 0, 40, 40, 40, 40, 40, 40, 
    40, 40, 999, 999, 999, 999, 999, 999, 999, 999, 0, 0, 999, 999, 999, 999, 
    999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 40, 
    40, 999, 999, 999, 999, 0, 0, 999, 999, 999, 999, 999, 999, 0, 0, 0, 0 ;

 fleafcn = 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 
    999, 999, 999, 999, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 
    65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 
    65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 
    65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65 ;

 fleafi = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0.8, 0.8, 0.75, 
    0.75, 0.425, 0.425, 0.85, 0.85, 0.75, 0.75, 0.425, 0.425, 0.75, 0.75, 
    0.425, 0.425, _, _, _, _, _, _, _, _, 0.85, 0.85, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, 0.75, 0.75, _, _, _, _, 0.8, 0.8, _, _, _, 
    _, _, _, 0.8, 0.8, 0.85, 0.85 ;

 flivewd = 0, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.5, 0.5, 0.1, 0, 0, 0, 
    0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 flnr = 0, 0.0509, 0.0466, 0.0546, 0.0461, 0.0515, 0.0716, 0.1007, 0.1007, 
    0.0517, 0.0943, 0.0943, 0.1365, 0.1365, 0.09, 0.1758, 0.1758, 0.293, 
    0.293, 0.4102, 0.4102, 0.4102, 0.4102, 0.4102, 0.4102, 0.4102, 0.4102, 
    0.4102, 0.4102, 0.4102, 0.4102, 0.4102, 0.4102, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.4102, 0.4102, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.4102, 0.4102, 0, 0, 0, 0, 0.293, 0.293, 0, 0, 0, 0, 0, 0, 0.293, 0.293, 
    0.4102, 0.4102 ;

 fm_droot = 0, 0.13, 0.15, 0.15, 0.13, 0.13, 0.1, 0.1, 0.13, 0.17, 0.17, 
    0.17, 0.2, 0.2, 0.2, 0.2, 0.2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 fm_dstem = 0, 0.45, 0.5, 0.5, 0.45, 0.45, 0.35, 0.35, 0.45, 0.55, 0.55, 
    0.55, 0.8, 0.8, 0.8, 0.8, 0.8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 fm_leaf = 0, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 
    0.8, 0.8, 0.8, 0.8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 fm_lroot = 0, 0.13, 0.15, 0.15, 0.13, 0.13, 0.1, 0.1, 0.13, 0.17, 0.17, 
    0.17, 0.2, 0.2, 0.2, 0.2, 0.2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 fm_lstem = 0, 0.45, 0.5, 0.5, 0.45, 0.45, 0.35, 0.35, 0.45, 0.55, 0.55, 
    0.55, 0.8, 0.8, 0.8, 0.8, 0.8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 fm_other = 0, 0.45, 0.5, 0.5, 0.45, 0.45, 0.35, 0.35, 0.45, 0.55, 0.55, 
    0.55, 0.8, 0.8, 0.8, 0.8, 0.8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 fm_root = 0, 0.13, 0.15, 0.15, 0.13, 0.13, 0.1, 0.1, 0.13, 0.17, 0.17, 0.17, 
    0.2, 0.2, 0.2, 0.2, 0.2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 fnitr = 0, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 
    50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 
    50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 
    50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 
    50, 50, 50, 50, 50, 50, 50, 50 ;

 fr_fcel = 0, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5 ;

 fr_flab = 0, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25 ;

 fr_flig = 0, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25 ;

 froot_leaf = 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2 ;

 frootcn = 1, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 
    42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 
    42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 
    42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 
    42, 42, 42, 42, 42, 42, 42, 42 ;

 frootcn_max = 1, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 
    52, 52, 52, 52, 52, 52, 52, 52, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 frootcn_min = 1, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 
    32, 32, 32, 32, 32, 32, 32, 32, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 froz_q10 = 1.5 ;

 fsr_pft = 0, 0.4, 0.43, 0.43, 0.4, 0.4, 0.4, 0.4, 0.4, 0.46, 0.46, 0.46, 
    0.6, 0.6, 0.6, 0.6, 0.6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 fstemcn = 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 
    999, 999, 999, 999, 120, 120, 100, 100, 100, 100, 130, 130, 100, 100, 
    100, 100, 100, 100, 100, 100, 999, 999, 999, 999, 999, 999, 999, 999, 
    130, 130, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 
    999, 999, 999, 999, 999, 999, 100, 100, 999, 999, 999, 999, 120, 120, 
    999, 999, 999, 999, 999, 999, 120, 120, 130, 130 ;

 fstor2tran = 0.5 ;

 fun_cn_flex_a = 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5 ;

 fun_cn_flex_b = 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 
    200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 
    200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 
    200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 
    200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 
    200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200 ;

 fun_cn_flex_c = 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 
    8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 
    8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 
    8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8 ;

 gddfunc_p1 = 4.8 ;

 gddfunc_p2 = 0.13 ;

 gddmin = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 50, 50, 50, 50, 
    50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 
    50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 
    50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 
    50, 50, 50, 50 ;

 graincn = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 50, 50, 50, 50, 
    50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 
    50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 
    50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 
    50, 50, 50, 50 ;

 grnfill = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0.65, 0.65, 
    0.6, 0.6, 0.4, 0.4, 0.7, 0.7, 0.6, 0.6, 0.4, 0.4, 0.6, 0.6, 0.4, 0.4, _, 
    _, _, _, _, _, _, _, 0.7, 0.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, 0.6, 0.6, _, _, _, _, 0.65, 0.65, _, _, _, _, _, _, 0.65, 
    0.65, 0.7, 0.7 ;

 grperc = 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 
    0.3, 0.3, 0.3, 0.3, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25 ;

 grpnow = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 highlatfact = 2 ;

 hybgdd = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 1700, 1700, 
    1700, 1700, 1700, 1700, 1900, 1900, 1700, 1700, 1700, 1700, 1700, 1700, 
    1700, 1700, _, _, _, _, _, _, _, _, 1700, 1700, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, 2100, 2100, _, _, _, _, 4300, 4300, _, _, 
    _, _, _, _, 1800, 1800, 2100, 2100 ;

 i_flnr = 0, 0.24, 0.24, 0.24, 0.18, 0.24, 0.18, 0.24, 0.24, 0.2, 0.2, 0.2, 
    0.28, 0.28, 0.28, 0.28, 0.28, 0.28, 0.28, 0.28, 0.28, 0.28, 0.28, 0.28, 
    0.28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0 ;

 i_vc = 0, 34.05, 34.05, 34.05, 1.99, 5.4, 6.35, 5.4, 5.4, 4.61, 4.61, 4.61, 
    23.74, 23.74, 23.74, 22.22, 22.22, 22.22, 22.22, 22.22, 22.22, 22.22, 
    22.22, 22.22, 22.22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 i_vca = 0, 6.32, 6.32, 6.32, 8.9, 5.73, 4.19, 5.73, 5.73, 14.71, 14.71, 
    14.71, 6.42, 6.42, 6.42, 4.71, 4.71, 4.71, 4.71, 4.71, 4.71, 4.71, 4.71, 
    4.71, 4.71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 i_vcad = 0, 6.32, 6.32, 6.32, 30.93, 5.73, 4.19, 5.73, 5.73, 14.71, 14.71, 
    14.71, 6.42, 6.42, 6.42, 4.71, 4.71, 4.71, 4.71, 4.71, 4.71, 4.71, 4.71, 
    4.71, 4.71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 irrigated = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 
    0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 
    0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 
    0, 1, 0, 1, 0, 1, 0, 1, 0, 1 ;

 k_frag = 0.00100050033358353 ;

 k_l1 = 1.20397280432594 ;

 k_l2 = 0.0725706928348355 ;

 k_l3 = 0.0140989243795016 ;

 k_m = 0.005 ;

 k_m_o2 = 0.02 ;

 k_m_unsat = 0.0005 ;

 k_mort = 0.3 ;

 k_nitr_max = 1.1574074e-06 ;

 k_s1 = 0.0725706928348355 ;

 k_s2 = 0.0140989243795016 ;

 k_s3 = 0.0014009809156281 ;

 k_s4 = 0.000100005000333347 ;

 kc_nonmyc = 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481, 0.000280893961280481, 
    0.000280893961280481, 0.000280893961280481 ;

 kmax =
  0, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07,
  0, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07,
  0, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07,
  0, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 
    1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07, 1e-07 ;

 kn_nonmyc = 0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042, 0.00328853498220042, 0.00328853498220042, 
    0.00328853498220042 ;

 kr_resorb = 0.00194149850039119, 0.00194149850039119, 0.00194149850039119, 
    9.6906331404746, 0.00194149850039119, 0.00194149850039119, 
    9.6906331404746, 9.6906331404746, 9.6906331404746, 0.00194149850039119, 
    9.6906331404746, 9.6906331404746, 9.6906331404746, 9.6906331404746, 
    9.6906331404746, 9.6906331404746, 9.6906331404746, 9.6906331404746, 
    9.6906331404746, 9.6906331404746, 9.6906331404746, 9.6906331404746, 
    9.6906331404746, 9.6906331404746, 9.6906331404746, 9.6906331404746, 
    9.6906331404746, 9.6906331404746, 9.6906331404746, 9.6906331404746, 
    9.6906331404746, 9.6906331404746, 9.6906331404746, 9.6906331404746, 
    9.6906331404746, 9.6906331404746, 9.6906331404746, 9.6906331404746, 
    9.6906331404746, 9.6906331404746, 9.6906331404746, 9.6906331404746, 
    9.6906331404746, 9.6906331404746, 9.6906331404746, 9.6906331404746, 
    9.6906331404746, 9.6906331404746, 9.6906331404746, 9.6906331404746, 
    9.6906331404746, 9.6906331404746, 9.6906331404746, 9.6906331404746, 
    9.6906331404746, 9.6906331404746, 9.6906331404746, 9.6906331404746, 
    9.6906331404746, 9.6906331404746, 9.6906331404746, 9.6906331404746, 
    9.6906331404746, 9.6906331404746, 9.6906331404746, 9.6906331404746, 
    9.6906331404746, 9.6906331404746, 9.6906331404746, 9.6906331404746, 
    9.6906331404746, 9.6906331404746, 9.6906331404746, 9.6906331404746, 
    9.6906331404746, 9.6906331404746, 9.6906331404746, 9.6906331404746, 
    9.6906331404746 ;

 krmax = 0, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 
    2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 
    2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 
    2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 
    2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 
    2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 
    2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 
    2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09, 2e-09 ;

 laimx = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 5, 5, 7, 7, 7, 7, 
    6, 6, 7, 7, 7, 7, 7, 7, 7, 7, _, _, _, _, _, _, _, _, 6, 6, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, 7, 7, _, _, _, _, 5, 5, _, _, 
    _, _, _, _, 5, 5, 6, 6 ;

 lake_decomp_fact = 9e-11 ;

 leaf_long = 0, 3, 6, 1, 1.5, 1.5, 1, 1, 1, 1.5, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 leafcn = 1, 35, 40, 25, 30, 30, 25, 25, 25, 30, 25, 25, 25, 25, 25, 25, 25, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25, 25, 25, 25, 25, 25, 25, 25 ;

 leafcn_max = 1, 45, 50, 35, 40, 40, 35, 35, 35, 40, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 leafcn_min = 1, 25, 30, 15, 20, 20, 15, 15, 15, 20, 15, 15, 15, 15, 15, 15, 
    15, 15, 15, 15, 15, 15, 15, 15, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 lf_fcel = 0, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5 ;

 lf_flab = 0, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25 ;

 lf_flig = 0, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25 ;

 lfemerg = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0.03, 0.03, 
    0.05, 0.05, 0.05, 0.05, 0.03, 0.03, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.05, _, _, _, _, _, _, _, _, 0.03, 0.03, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, 0.05, 0.05, _, _, _, _, 0.03, 0.03, _, _, 
    _, _, _, _, 0.03, 0.03, 0.03, 0.03 ;

 lflitcn = 1, 70, 80, 50, 60, 60, 50, 50, 50, 60, 50, 50, 50, 50, 50, 50, 50, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 
    25, 25, 25, 25, 25, 25, 25, 25 ;

 lfr_cn = 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 
    0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0 ;

 livewdcn = 1, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 0, 0, 0, 0, 0, 50, 
    50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 
    50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 
    50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 
    50, 50, 50, 50, 50, 50, 50 ;

 livewdcn_max = 1, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 0, 0, 0, 0, 0, 
    60, 60, 60, 60, 60, 60, 60, 60, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 livewdcn_min = 1, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 0, 0, 0, 0, 0, 
    40, 40, 40, 40, 40, 40, 40, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 lmr_intercept_atkin = 0, 1.4995, 1.4995, 1.4995, 1.756, 1.756, 1.756, 1.756, 
    1.756, 2.0749, 2.0749, 2.0749, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 
    2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 
    2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 
    2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 
    2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 
    2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 
    2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 
    2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956, 2.1956 ;

 lwtop_ann = 0.7 ;

 max_NH_planting_date = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    615, 615, 615, 615, 1130, 1130, 615, 615, 615, 615, 1130, 1130, 615, 615, 
    1130, 1130, _, _, _, _, _, _, _, _, 531, 531, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, 228, 228, _, _, _, _, 331, 331, _, _, _, _, _, 
    _, 415, 415, 701, 701 ;

 max_SH_planting_date = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    1215, 1215, 1215, 1215, 530, 530, 1215, 1215, 1215, 1215, 530, 530, 1215, 
    1215, 530, 530, _, _, _, _, _, _, _, _, 1130, 1130, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, 1231, 1231, _, _, _, _, 1031, 1031, _, 
    _, _, _, _, _, 1015, 1015, 1231, 1231 ;

 max_altdepth_cryoturbation = 2 ;

 max_altmultiplier_cryoturb = 3 ;

 maxpsi_hr = -0.03 ;

 mbbopt = 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 4, 9, 9, 4, 4, 9, 9, 9, 
    9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 
    9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 4, 4, 9, 
    9, 9, 9, 9, 9, 4, 4, 9, 9 ;

 me_herb = 0.2 ;

 me_woody = 0.3 ;

 mergetoclmpft = _, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 
    17, 18, 19, 20, 21, 22, 23, 24, 19, 20, 21, 22, 19, 20, 21, 22, 15, 16, 
    15, 16, 15, 16, 15, 16, 41, 42, 15, 16, 15, 16, 15, 16, 15, 16, 15, 16, 
    15, 16, 15, 16, 15, 16, 15, 16, 61, 62, 15, 16, 15, 16, 67, 68, 15, 16, 
    15, 16, 15, 16, 75, 76, 77, 78 ;

 min_NH_planting_date = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    401, 401, 401, 401, 901, 901, 501, 501, 401, 401, 901, 901, 401, 401, 
    901, 901, _, _, _, _, _, _, _, _, 401, 401, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, 101, 101, _, _, _, _, 101, 101, _, _, _, _, _, _, 
    320, 320, 415, 415 ;

 min_SH_planting_date = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    1001, 1001, 1001, 1001, 301, 301, 1101, 1101, 1001, 1001, 301, 301, 1001, 
    1001, 301, 301, _, _, _, _, _, _, _, _, 901, 901, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, 1015, 1015, _, _, _, _, 801, 801, _, _, _, 
    _, _, _, 920, 920, 1015, 1015 ;

 min_planting_temp = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    279.15, 279.15, 272.15, 272.15, 278.15, 278.15, 279.15, 279.15, 272.15, 
    272.15, 278.15, 278.15, 272.15, 272.15, 278.15, 278.15, _, _, _, _, _, _, 
    _, _, 283.15, 283.15, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, 283.15, 283.15, _, _, _, _, 283.15, 283.15, _, _, _, _, _, _, 283.15, 
    283.15, 283.15, 283.15 ;

 minfuel = 100 ;

 mino2lim = 0.2 ;

 minpsi_hr = -10 ;

 mxmat = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 165, 165, 150, 
    150, 265, 265, 150, 150, 150, 150, 265, 265, 150, 150, 265, 265, _, _, _, 
    _, _, _, _, _, 160, 160, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, 150, 150, _, _, _, _, 300, 300, _, _, _, _, _, _, 160, 160, 150, 150 ;

 mxtmp = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 30, 30, 26, 26, 
    26, 26, 30, 30, 26, 26, 26, 26, 26, 26, 26, 26, _, _, _, _, _, _, _, _, 
    30, 30, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 30, 30, _, 
    _, _, _, 30, 30, _, _, _, _, _, _, 30, 30, 30, 30 ;

 ndays_off = 15 ;

 ndays_on = 30 ;

 nfr_cn = 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0 ;

 nongrassporosratio = 0.33 ;

 organic_max = 130 ;

 oxinhib = 400 ;

 pHmax = 9 ;

 pHmin = 2.2 ;

 pconv = 0, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.8, 0.8, 0.8, 1, 1, 1, 
    1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 perecm = 1, 1, 1, 1, 0, 0, 0, 0.5, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 pftname =
  "not_vegetated                           ",
  "needleleaf_evergreen_temperate_tree     ",
  "needleleaf_evergreen_boreal_tree        ",
  "needleleaf_deciduous_boreal_tree        ",
  "broadleaf_evergreen_tropical_tree       ",
  "broadleaf_evergreen_temperate_tree      ",
  "broadleaf_deciduous_tropical_tree       ",
  "broadleaf_deciduous_temperate_tree      ",
  "broadleaf_deciduous_boreal_tree         ",
  "broadleaf_evergreen_shrub               ",
  "broadleaf_deciduous_temperate_shrub     ",
  "broadleaf_deciduous_boreal_shrub        ",
  "c3_arctic_grass                         ",
  "c3_non-arctic_grass                     ",
  "c4_grass                                ",
  "c3_crop                                 ",
  "c3_irrigated                            ",
  "temperate_corn                          ",
  "irrigated_temperate_corn                ",
  "spring_wheat                            ",
  "irrigated_spring_wheat                  ",
  "winter_wheat                            ",
  "irrigated_winter_wheat                  ",
  "temperate_soybean                       ",
  "irrigated_temperate_soybean             ",
  "barley                                  ",
  "irrigated_barley                        ",
  "winter_barley                           ",
  "irrigated_winter_barley                 ",
  "rye                                     ",
  "irrigated_rye                           ",
  "winter_rye                              ",
  "irrigated_winter_rye                    ",
  "cassava                                 ",
  "irrigated_cassava                       ",
  "citrus                                  ",
  "irrigated_citrus                        ",
  "cocoa                                   ",
  "irrigated_cocoa                         ",
  "coffee                                  ",
  "irrigated_coffee                        ",
  "cotton                                  ",
  "irrigated_cotton                        ",
  "datepalm                                ",
  "irrigated_datepalm                      ",
  "foddergrass                             ",
  "irrigated_foddergrass                   ",
  "grapes                                  ",
  "irrigated_grapes                        ",
  "groundnuts                              ",
  "irrigated_groundnuts                    ",
  "millet                                  ",
  "irrigated_millet                        ",
  "oilpalm                                 ",
  "irrigated_oilpalm                       ",
  "potatoes                                ",
  "irrigated_potatoes                      ",
  "pulses                                  ",
  "irrigated_pulses                        ",
  "rapeseed                                ",
  "irrigated_rapeseed                      ",
  "rice                                    ",
  "irrigated_rice                          ",
  "sorghum                                 ",
  "irrigated_sorghum                       ",
  "sugarbeet                               ",
  "irrigated_sugarbeet                     ",
  "sugarcane                               ",
  "irrigated_sugarcane                     ",
  "sunflower                               ",
  "irrigated_sunflower                     ",
  "miscanthus                              ",
  "irrigated_miscanthus                    ",
  "switchgrass                             ",
  "irrigated_switchgrass                   ",
  "tropical_corn                           ",
  "irrigated_tropical_corn                 ",
  "tropical_soybean                        ",
  "irrigated_tropical_soybean              " ;

 pftnum = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78 ;

 pftpar20 = _, 15, 15, 15, 15, 15, 15, 15, 15, 5, 5, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 pftpar28 = _, -2, -32.5, _, 15.5, 3, 15.5, -17, -1000, _, -17, -1000, -1000, 
    -17, 15.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 pftpar29 = _, 22, -2, -2, _, 18.8, _, 15.5, -2, _, _, -2, -17, 15.5, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 pftpar30 = 0, 900, 600, 350, 0, 1200, 0, 1200, 350, 0, 1200, 350, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 pftpar31 = _, _, 23, 23, _, _, _, _, 23, _, _, 23, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _ ;

 planting_temp = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 283.15, 
    283.15, 280.15, 280.15, _, _, 286.15, 286.15, 280.15, 280.15, _, _, 
    280.15, 280.15, _, _, _, _, _, _, _, _, _, _, 294.15, 294.15, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, 294.15, 294.15, _, _, _, _, 
    294.15, 294.15, _, _, _, _, _, _, 294.15, 294.15, 294.15, 294.15 ;

 porosmin = 0.05 ;

 pprod10 = 0, 0.3, 0.3, 0.3, 0.4, 0.3, 0.4, 0.3, 0.3, 0.2, 0.2, 0.2, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 pprod100 = 0, 0.1, 0.1, 0.1, 0, 0.1, 0, 0.1, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 pprodharv10 = _, 0.75, 0.75, 0.75, 1, 0.75, 1, 0.75, 0.75, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 psi50 =
  0, -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000,
  0, -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000,
  0, -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000,
  0, -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000, -200000, -200000, 
    -200000, -200000, -200000, -200000, -200000, -200000 ;

 psi_soil_ref = 0, -50000, -50000, -50000, -50000, -50000, -50000, -50000, 
    -50000, -50000, -50000, -50000, -50000, -50000, -50000, -50000, -50000, 
    -50000, -50000, -50000, -50000, -50000, -50000, -50000, -50000, -50000, 
    -50000, -50000, -50000, -50000, -50000, -50000, -50000, -50000, -50000, 
    -50000, -50000, -50000, -50000, -50000, -50000, -50000, -50000, -50000, 
    -50000, -50000, -50000, -50000, -50000, -50000, -50000, -50000, -50000, 
    -50000, -50000, -50000, -50000, -50000, -50000, -50000, -50000, -50000, 
    -50000, -50000, -50000, -50000, -50000, -50000, -50000, -50000, -50000, 
    -50000, -50000, -50000, -50000, -50000, -50000, -50000, -50000 ;

 q10_ch4oxid = 1.9 ;

 q10_hr = 1.5 ;

 q10_mr = 1.5 ;

 q10ch4 = 1.33 ;

 q10ch4base = 295 ;

 q10lakebase = 298 ;

 qflxlagd = 30 ;

 r_mort = 0.02 ;

 rc_npool = 10 ;

 redoxlag = 30 ;

 redoxlag_vertical = 0 ;

 rf_cwdl2_bgc = 0 ;

 rf_cwdl3_bgc = 0 ;

 rf_l1s1 = 0.39 ;

 rf_l1s1_bgc = 0.55 ;

 rf_l2s1_bgc = 0.5 ;

 rf_l2s2 = 0.55 ;

 rf_l3s2_bgc = 0.5 ;

 rf_l3s3 = 0.29 ;

 rf_s1s2 = 0.28 ;

 rf_s2s1_bgc = 0.55 ;

 rf_s2s3 = 0.46 ;

 rf_s2s3_bgc = 0.55 ;

 rf_s3s1_bgc = 0.55 ;

 rf_s3s4 = 0.55 ;

 rholnir = 0, 0.35, 0.35, 0.35, 0.45, 0.45, 0.45, 0.45, 0.45, 0.35, 0.45, 
    0.45, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 
    0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 
    0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.58, 0.58, 0.35, 0.35, 0.35, 0.35, 
    0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 0.35, 
    0.35, 0.35, 0.58, 0.58, 0.35, 0.35, 0.35, 0.35, 0.58, 0.58, 0.35, 0.35, 
    0.35, 0.35, 0.35, 0.35, 0.58, 0.58, 0.58, 0.58 ;

 rholvis = 0, 0.07, 0.07, 0.07, 0.1, 0.1, 0.1, 0.1, 0.1, 0.07, 0.1, 0.1, 
    0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 
    0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 
    0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 
    0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 
    0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 
    0.11, 0.11, 0.11, 0.11, 0.11, 0.11, 0.11 ;

 rhosnir = 0, 0.39, 0.39, 0.39, 0.39, 0.39, 0.39, 0.39, 0.39, 0.39, 0.39, 
    0.39, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 
    0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 
    0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 
    0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 
    0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 
    0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53, 0.53 ;

 rhosvis = 0, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 
    0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 
    0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 
    0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 
    0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 
    0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31, 0.31 ;

 rij_kro_a = 1.5e-10 ;

 rij_kro_alpha = 1.26 ;

 rij_kro_beta = 0.6 ;

 rij_kro_delta = 0.85 ;

 rij_kro_gamma = 0.6 ;

 rob = 3 ;

 root_dmx = 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 
    999, 999, 999, 999, 1.20000004768372, 1.20000004768372, 
    0.899999976158142, 0.899999976158142, 0.899999976158142, 
    0.899999976158142, 1.60000002384186, 1.60000002384186, 1.60000002384186, 
    1.60000002384186, 1.60000002384186, 1.60000002384186, 1.60000002384186, 
    1.60000002384186, 1.60000002384186, 1.60000002384186, 1.60000002384186, 
    1.60000002384186, 1.60000002384186, 1.60000002384186, 1.60000002384186, 
    1.60000002384186, 1.60000002384186, 1.60000002384186, 1.60000002384186, 
    1.60000002384186, 1.60000002384186, 1.60000002384186, 1.60000002384186, 
    1.60000002384186, 1.60000002384186, 1.60000002384186, 1.60000002384186, 
    1.60000002384186, 1.60000002384186, 1.60000002384186, 1.60000002384186, 
    1.60000002384186, 1.60000002384186, 1.60000002384186, 1.60000002384186, 
    1.60000002384186, 1.60000002384186, 1.60000002384186, 1.60000002384186, 
    1.60000002384186, 1.60000002384186, 1.60000002384186, 1.60000002384186, 
    1.60000002384186, 1.60000002384186, 1.60000002384186, 1.60000002384186, 
    1.60000002384186, 1.60000002384186, 1.60000002384186, 1.60000002384186, 
    1.60000002384186, 1.60000002384186, 1.60000002384186, 1.60000002384186, 
    1.60000002384186 ;

 roota_par = 0, 7, 7, 7, 7, 7, 6, 6, 6, 7, 7, 7, 11, 11, 11, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6 ;

 rootb_par = 0, 2, 2, 2, 1, 1, 2, 2, 2, 1.5, 1.5, 1.5, 2, 2, 2, 3, 3, 3, 3, 
    3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 
    3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 
    3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3 ;

 rootlitfrac = 0.5 ;

 s_fix = -14.456888485725, -14.456888485725, -14.456888485725, 
    -14.456888485725, -14.456888485725, -14.456888485725, -14.456888485725, 
    -14.456888485725, -14.456888485725, -14.456888485725, -14.456888485725, 
    -14.456888485725, -14.456888485725, -14.456888485725, -14.456888485725, 
    -14.456888485725, -14.456888485725, -14.456888485725, -14.456888485725, 
    -14.456888485725, -14.456888485725, -14.456888485725, -14.456888485725, 
    -14.456888485725, -14.456888485725, -14.456888485725, -14.456888485725, 
    -14.456888485725, -14.456888485725, -14.456888485725, -14.456888485725, 
    -14.456888485725, -14.456888485725, -14.456888485725, -14.456888485725, 
    -14.456888485725, -14.456888485725, -14.456888485725, -14.456888485725, 
    -14.456888485725, -14.456888485725, -14.456888485725, -14.456888485725, 
    -14.456888485725, -14.456888485725, -14.456888485725, -14.456888485725, 
    -14.456888485725, -14.456888485725, -14.456888485725, -14.456888485725, 
    -14.456888485725, -14.456888485725, -14.456888485725, -14.456888485725, 
    -14.456888485725, -14.456888485725, -14.456888485725, -14.456888485725, 
    -14.456888485725, -14.456888485725, -14.456888485725, -14.456888485725, 
    -14.456888485725, -14.456888485725, -14.456888485725, -14.456888485725, 
    -14.456888485725, -14.456888485725, -14.456888485725, -14.456888485725, 
    -14.456888485725, -14.456888485725, -14.456888485725, -14.456888485725, 
    -14.456888485725, -14.456888485725, -14.456888485725, -14.456888485725 ;

 s_flnr = 0, -0.22, -0.22, -0.22, -0.38, -0.22, -0.38, -0.22, -0.22, -0.01, 
    -0.01, -0.01, -0.03, -0.03, -0.03, -0.03, -0.03, -0.03, -0.03, -0.03, 
    -0.03, -0.03, -0.03, -0.03, -0.03, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 s_vc = 0, 9.71, 9.71, 9.71, 10.71, 30.38, 25.88, 30.38, 30.38, 30.2, 30.2, 
    30.2, 28.17, 28.17, 28.17, 41.27, 41.27, 41.27, 41.27, 41.27, 41.27, 
    41.27, 41.27, 41.27, 41.27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 s_vca = 0, 18.15, 18.15, 18.15, 9.3, 29.81, 26.19, 29.81, 29.81, 23.15, 
    23.15, 23.15, 40.96, 40.96, 40.96, 59.23, 59.23, 59.23, 59.23, 59.23, 
    59.23, 59.23, 59.23, 59.23, 59.23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 s_vcad = 0, 18.15, 18.15, 18.15, 5.5, 29.81, 26.19, 29.81, 29.81, 23.15, 
    23.15, 23.15, 40.96, 40.96, 40.96, 59.23, 59.23, 59.23, 59.23, 59.23, 
    59.23, 59.23, 59.23, 59.23, 59.23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 satpow = 2 ;

 scale_factor_aere = 1 ;

 scale_factor_gasdiff = 1 ;

 scale_factor_liqdiff = 1 ;

 season_decid = 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 segment =
  "sunlit                                  ",
  "shaded                                  ",
  "xylem                                   ",
  "root                                    " ;

 sf_minn = 0.1 ;

 sf_no3 = 1 ;

 shape_fluxprof_param1 = 10000000000 ;

 slatop = 0, 0.01, 0.008, 0.024, 0.012, 0.012, 0.03, 0.03, 0.03, 0.012, 0.03, 
    0.03, 0.03, 0.03, 0.03, 0.03, 0.03, 0.05, 0.05, 0.07, 0.07, 0.07, 0.07, 
    0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.07, 0.07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.07, 0.07, 0, 0, 0, 0, 0.05, 0.05, 0, 0, 0, 0, 0, 0, 0.05, 0.05, 
    0.07, 0.07 ;

 smp_crit = -240000 ;

 smpsc = 0, -255000, -255000, -255000, -255000, -255000, -224000, -224000, 
    -224000, -428000, -428000, -428000, -275000, -275000, -275000, -275000, 
    -275000, -275000, -275000, -275000, -275000, -275000, -275000, -275000, 
    -275000, -275000, -275000, -275000, -275000, -275000, -275000, -275000, 
    -275000, -275000, -275000, -275000, -275000, -275000, -275000, -275000, 
    -275000, -275000, -275000, -275000, -275000, -275000, -275000, -275000, 
    -275000, -275000, -275000, -275000, -275000, -275000, -275000, -275000, 
    -275000, -275000, -275000, -275000, -275000, -275000, -275000, -275000, 
    -275000, -275000, -275000, -275000, -275000, -275000, -275000, -275000, 
    -275000, -275000, -275000, -275000, -275000, -275000, -275000 ;

 smpso = 0, -66000, -66000, -66000, -66000, -66000, -35000, -35000, -35000, 
    -83000, -83000, -83000, -74000, -74000, -74000, -74000, -74000, -74000, 
    -74000, -74000, -74000, -74000, -74000, -74000, -74000, -74000, -74000, 
    -74000, -74000, -74000, -74000, -74000, -74000, -74000, -74000, -74000, 
    -74000, -74000, -74000, -74000, -74000, -74000, -74000, -74000, -74000, 
    -74000, -74000, -74000, -74000, -74000, -74000, -74000, -74000, -74000, 
    -74000, -74000, -74000, -74000, -74000, -74000, -74000, -74000, -74000, 
    -74000, -74000, -74000, -74000, -74000, -74000, -74000, -74000, -74000, 
    -74000, -74000, -74000, -74000, -74000, -74000, -74000 ;

 soilpsi_off = -2 ;

 soilpsi_on = -2 ;

 som_diffus = 3.171e-12 ;

 stem_leaf = 0, -1, -1, -1, -1, -1, -1, -1, -1, 0.2, 0.2, 0.2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 stress_decid = 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 surface_tension_water = 0.073 ;

 tau_cwd = 3.3333333333333 ;

 tau_l1 = 0.054054054054 ;

 tau_l2_l3 = 0.204081632653061 ;

 tau_s1 = 0.136986301369863 ;

 tau_s2 = 5 ;

 tau_s3 = 222.222222222222 ;

 taulnir = 0, 0.1, 0.1, 0.1, 0.25, 0.25, 0.25, 0.25, 0.25, 0.1, 0.25, 0.25, 
    0.34, 0.34, 0.34, 0.34, 0.34, 0.34, 0.34, 0.34, 0.34, 0.34, 0.34, 0.34, 
    0.34, 0.34, 0.34, 0.34, 0.34, 0.34, 0.34, 0.34, 0.34, 0.34, 0.34, 0.34, 
    0.34, 0.34, 0.34, 0.34, 0.34, 0.25, 0.25, 0.34, 0.34, 0.34, 0.34, 0.34, 
    0.34, 0.34, 0.34, 0.34, 0.34, 0.34, 0.34, 0.34, 0.34, 0.34, 0.34, 0.34, 
    0.34, 0.25, 0.25, 0.34, 0.34, 0.34, 0.34, 0.25, 0.25, 0.34, 0.34, 0.34, 
    0.34, 0.34, 0.34, 0.25, 0.25, 0.25, 0.25 ;

 taulvis = 0, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.07, 0.07, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 0.05, 
    0.05, 0.05, 0.07, 0.07, 0.05, 0.05, 0.05, 0.05, 0.07, 0.07, 0.05, 0.05, 
    0.05, 0.05, 0.05, 0.05, 0.07, 0.07, 0.07, 0.07 ;

 tausnir = 0, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 
    0.001, 0.001, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 
    0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25, 0.25 ;

 tausvis = 0, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 
    0.001, 0.001, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 
    0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 
    0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 
    0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 
    0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 
    0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12 ;

 unsat_aere_ratio = 0.166666666666667 ;

 vgc_max = 0.15 ;

 vmax_ch4_oxid = 1.25e-05 ;

 vmax_oxid_unsat = 1.25e-06 ;

 wcf = 0.4 ;

 woody = 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0 ;

 xl = 0, 0.01, 0.01, 0.01, 0.1, 0.1, 0.01, 0.25, 0.25, 0.01, 0.25, 0.25, 
    -0.3, -0.3, -0.3, -0.3, -0.3, -0.5, -0.5, 0.65, 0.65, 0.65, 0.65, -0.5, 
    -0.5, 0.65, 0.65, 0.65, 0.65, 0.65, 0.65, 0.65, 0.65, 0, 0, 0, 0, 0, 0, 
    0, 0, -0.5, -0.5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.65, 0.65, 0, 0, 0, 0, -0.5, -0.5, 0, 0, 0, 0, 0, 0, -0.5, -0.5, -0.5, 
    -0.5 ;

 z0mr = 0, 0.055, 0.055, 0.055, 0.075, 0.075, 0.055, 0.055, 0.055, 0.12, 
    0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 
    0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 
    0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 
    0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 
    0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 
    0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12, 0.12 ;

 ztopmx = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2.5, 2.5, 1.2, 
    1.2, 1.2, 1.2, 0.75, 0.75, 1.2, 1.2, 1.2, 1.2, 1.2, 1.2, 1.2, 1.2, _, _, 
    _, _, _, _, _, _, 1.5, 1.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, 1.8, 1.8, _, _, _, _, 4, 4, _, _, _, _, _, _, 2.5, 2.5, 1, 1 ;

 rootprof_beta =
  0, 0.976, 0.943, 0.943, 0.993, 0.966, 0.993, 0.966, 0.943, 0.964, 0.964, 
    0.914, 0.914, 0.943, 0.943, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 
    0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 
    0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 
    0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 
    0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 
    0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 
    0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961,
  0, 0.976, 0.943, 0.943, 0.962, 0.966, 0.961, 0.966, 0.943, 0.964, 0.964, 
    0.914, 0.914, 0.943, 0.943, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 
    0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 
    0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 
    0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 
    0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 
    0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 
    0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961, 0.961 ;

 wood_density = 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 
    0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _ ;

 BB_slope = 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 
    8, 8, 8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _ ;

 alpha_stem = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _ ;

 leaf_stor_priority = 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 
    0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _ ;

 max_dbh = 68, 1.5, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 
    68, 68, 68, 68, 68, 68, 68, 68, 68, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 cushion = 1.2, 1.2, 1.2, 1.2, 1.2, 1.2, 1.2, 1.2, 1.2, 1.2, 1.2, 1.2, 1.2, 
    1.2, 1.2, 1.2, 1.2, 1.2, 1.2, 1.2, 1.2, 1.2, 1.2, 1.2, 1.2, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _ ;

 hgt_min = 1.25, 1.25, 1.25, 1.25, 1.25, 1.25, 1.25, 1.25, 1.25, 1.25, 1.25, 
    1.25, 1.25, 1.25, 1.25, 1.25, 1.25, 1.25, 1.25, 1.25, 1.25, 1.25, 1.25, 
    1.25, 1.25, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _ ;

 freezetol = 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 
    1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 
    1000, 1000, 1000, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _ ;

 resp_drought_response = 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _ ;

 leafwatermax = 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 
    0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _ ;

 rootresist = 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 
    200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _ ;

 soilbeta = 2000, 2000, 2000, 2000, 2000, 2000, 2000, 2000, 2000, 2000, 2000, 
    2000, 2000, 2000, 2000, 2000, 2000, 2000, 2000, 2000, 2000, 2000, 2000, 
    2000, 2000, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _ ;

 crown = 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _ ;

 bark_scaler = 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 
    0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 0.07, 
    0.07, 0.07, 0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _ ;

 crown_kill = 0.775, 0.775, 0.775, 0.775, 0.775, 0.775, 0.775, 0.775, 0.775, 
    0.775, 0.775, 0.775, 0.775, 0.775, 0.775, 0.775, 0.775, 0.775, 0.775, 
    0.775, 0.775, 0.775, 0.775, 0.775, 0.775, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 initd = 0.08, 0.06, 0.08, 0.08, 0.08, 0.08, 0.08, 0.08, 0.08, 0.08, 0.08, 
    0.08, 0.08, 0.08, 0.08, 0.08, 0.08, 0.08, 0.08, 0.08, 0.08, 0.08, 0.08, 
    0.08, 0.08, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _ ;

 sd_mort = 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 
    0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 
    0.98, 0.98, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _ ;

 seed_rain = 0.28, 0.28, 0.28, 0.28, 0.28, 0.28, 0.28, 0.28, 0.28, 0.28, 
    0.28, 0.28, 0.28, 0.28, 0.28, 0.28, 0.28, 0.28, 0.28, 0.28, 0.28, 0.28, 
    0.28, 0.28, 0.28, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _ ;

 bb_slope = 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _ ;

 root_long = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _ ;

 seed_alloc = 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 
    0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _ ;

 clone_alloc = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _ ;

 sapwood_ratio = 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 
    0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 
    0.001, 0.001, 0.001, 0.001, 0.001, 0.001, 0.001, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 grass_spread = 0.18 ;

 comp_excln = 0.1 ;

 stress_mort = 0.6 ;

 dispersal = 0.5 ;

 gr_perc = 0.2 ;

 maxspread = 0.3 ;

 minspread = 0.18 ;

 init_litter = 0.05 ;

 nfires = 15 ;

 understorey_death = 0.55983 ;

 profile_tol = 0.7 ;

 ag_biomass = 0.6 ;

 alpha_FMC = 0.00508, 0.001, 0.00028, 0.0008, 0.0004, 999 ;

 SAV = 66, 13, 3.58, 0.98, 0.2, 66 ;

 FBD = 4, 15.4, 16.8, 19.6, 999, 4 ;

 max_decomp = 1, 0.052, 0.016, 0.01, 0.0152, 999 ;

 min_moisture = 0.18, 0.15, 0.12, 0, 0, 0.18 ;

 mid_moisture = 0.73, 0.6, 0.51, 0.38, 0, 0.73 ;

 low_moisture_C = 1.1, 1.1, 2, 1.09, 0.98, 1.1 ;

 low_moisture_S = 0.62, 0.67, 0.72, 0.85, 0, 0.62 ;

 mid_moisture_C = 2.45, 2, 1.47, 1.06, 1, 2.45 ;

 mid_moisture_S = 2.45, 2, 1.47, 1.06, 0.8, 2.45 ;

 CWD_frac = 0.045, 0.075, 0.21, 0.67 ;

 fdi_a = 17.27 ;

 fdi_b = 237.7 ;

 fdi_alpha = 0.00037 ;

 miner_total = 0.055 ;

 fuel_energy = 18000 ;

 part_dens = 513 ;

 miner_damp = 0.055 ;

 max_durat = 240 ;

 durat_slope = -11.06 ;

 alpha_SH = 0.2 ;
}
